library verilog;
use verilog.vl_types.all;
entity alt_vipitc130_IS2Vid_calculate_mode is
    port(
        trs             : in     vl_logic_vector(3 downto 0);
        is_interlaced   : in     vl_logic;
        is_serial_output: in     vl_logic;
        is_sample_count_f0: in     vl_logic_vector(15 downto 0);
        is_line_count_f0: in     vl_logic_vector(15 downto 0);
        is_sample_count_f1: in     vl_logic_vector(15 downto 0);
        is_line_count_f1: in     vl_logic_vector(15 downto 0);
        is_h_front_porch: in     vl_logic_vector(15 downto 0);
        is_h_sync_length: in     vl_logic_vector(15 downto 0);
        is_h_blank      : in     vl_logic_vector(15 downto 0);
        is_v_front_porch: in     vl_logic_vector(15 downto 0);
        is_v_sync_length: in     vl_logic_vector(15 downto 0);
        is_v_blank      : in     vl_logic_vector(15 downto 0);
        is_v1_front_porch: in     vl_logic_vector(15 downto 0);
        is_v1_sync_length: in     vl_logic_vector(15 downto 0);
        is_v1_blank     : in     vl_logic_vector(15 downto 0);
        is_ap_line      : in     vl_logic_vector(15 downto 0);
        is_v1_rising_edge: in     vl_logic_vector(15 downto 0);
        is_f_rising_edge: in     vl_logic_vector(15 downto 0);
        is_f_falling_edge: in     vl_logic_vector(15 downto 0);
        is_anc_line     : in     vl_logic_vector(15 downto 0);
        is_v1_anc_line  : in     vl_logic_vector(15 downto 0);
        interlaced_nxt  : out    vl_logic;
        serial_output_nxt: out    vl_logic;
        h_total_minus_one_nxt: out    vl_logic_vector(15 downto 0);
        v_total_minus_one_nxt: out    vl_logic_vector(15 downto 0);
        ap_line_nxt     : out    vl_logic_vector(15 downto 0);
        ap_line_end_nxt : out    vl_logic_vector(15 downto 0);
        h_blank_nxt     : out    vl_logic_vector(15 downto 0);
        sav_nxt         : out    vl_logic_vector(15 downto 0);
        h_sync_start_nxt: out    vl_logic_vector(15 downto 0);
        h_sync_end_nxt  : out    vl_logic_vector(15 downto 0);
        f2_v_start_nxt  : out    vl_logic_vector(15 downto 0);
        f1_v_start_nxt  : out    vl_logic_vector(15 downto 0);
        f1_v_end_nxt    : out    vl_logic_vector(15 downto 0);
        f2_v_sync_start_nxt: out    vl_logic_vector(15 downto 0);
        f2_v_sync_end_nxt: out    vl_logic_vector(15 downto 0);
        f1_v_sync_start_nxt: out    vl_logic_vector(15 downto 0);
        f1_v_sync_end_nxt: out    vl_logic_vector(15 downto 0);
        f_rising_edge_nxt: out    vl_logic_vector(15 downto 0);
        f_falling_edge_nxt: out    vl_logic_vector(15 downto 0);
        total_line_count_f0_nxt: out    vl_logic_vector(12 downto 0);
        total_line_count_f1_nxt: out    vl_logic_vector(12 downto 0);
        f2_anc_v_start_nxt: out    vl_logic_vector(15 downto 0);
        f1_anc_v_start_nxt: out    vl_logic_vector(15 downto 0)
    );
end alt_vipitc130_IS2Vid_calculate_mode;
