library verilog;
use verilog.vl_types.all;
entity FFXII_LB_Cursor is
    generic(
        Y0X0            : integer := 0;
        Y0X1            : integer := 1;
        Y0X2            : integer := 2;
        Y0X3            : integer := 3;
        Y0X4            : integer := 4;
        Y0X5            : integer := 5;
        Y0X6            : integer := 6;
        Y0X7            : integer := 7;
        Y0X8            : integer := 8;
        Y0X9            : integer := 9;
        Y0X10           : integer := 10;
        Y0X11           : integer := 11;
        Y0X12           : integer := 12;
        Y0X13           : integer := 13;
        Y0X14           : integer := 14;
        Y0X15           : integer := 15;
        Y0X16           : integer := 16;
        Y0X17           : integer := 17;
        Y0X18           : integer := 18;
        Y0X19           : integer := 19;
        Y0X20           : integer := 20;
        Y0X21           : integer := 21;
        Y0X22           : integer := 22;
        Y0X23           : integer := 23;
        Y0X24           : integer := 24;
        Y0X25           : integer := 25;
        Y0X26           : integer := 26;
        Y0X27           : integer := 27;
        Y0X28           : integer := 28;
        Y1X1            : integer := 1025;
        Y1X2            : integer := 1026;
        Y1X3            : integer := 1027;
        Y1X4            : integer := 1028;
        Y1X5            : integer := 1029;
        Y1X6            : integer := 1030;
        Y1X7            : integer := 1031;
        Y1X8            : integer := 1032;
        Y1X9            : integer := 1033;
        Y1X10           : integer := 1034;
        Y1X11           : integer := 1035;
        Y1X12           : integer := 1036;
        Y1X13           : integer := 1037;
        Y1X14           : integer := 1038;
        Y1X15           : integer := 1039;
        Y1X16           : integer := 1040;
        Y1X17           : integer := 1041;
        Y1X18           : integer := 1042;
        Y1X19           : integer := 1043;
        Y1X20           : integer := 1044;
        Y1X21           : integer := 1045;
        Y1X22           : integer := 1046;
        Y1X23           : integer := 1047;
        Y1X24           : integer := 1048;
        Y1X25           : integer := 1049;
        Y1X26           : integer := 1050;
        Y1X27           : integer := 1051;
        Y1X28           : integer := 1052;
        Y2X1            : integer := 2049;
        Y2X2            : integer := 2050;
        Y2X3            : integer := 2051;
        Y2X4            : integer := 2052;
        Y2X5            : integer := 2053;
        Y2X6            : integer := 2054;
        Y2X7            : integer := 2055;
        Y2X8            : integer := 2056;
        Y2X9            : integer := 2057;
        Y2X10           : integer := 2058;
        Y2X11           : integer := 2059;
        Y2X12           : integer := 2060;
        Y2X13           : integer := 2061;
        Y2X14           : integer := 2062;
        Y2X15           : integer := 2063;
        Y2X16           : integer := 2064;
        Y2X17           : integer := 2065;
        Y2X18           : integer := 2066;
        Y2X19           : integer := 2067;
        Y2X20           : integer := 2068;
        Y2X21           : integer := 2069;
        Y2X22           : integer := 2070;
        Y2X23           : integer := 2071;
        Y2X24           : integer := 2072;
        Y2X25           : integer := 2073;
        Y2X26           : integer := 2074;
        Y2X27           : integer := 2075;
        Y2X28           : integer := 2076;
        Y3X1            : integer := 3073;
        Y3X2            : integer := 3074;
        Y3X3            : integer := 3075;
        Y3X4            : integer := 3076;
        Y3X5            : integer := 3077;
        Y3X6            : integer := 3078;
        Y3X7            : integer := 3079;
        Y3X8            : integer := 3080;
        Y3X9            : integer := 3081;
        Y3X10           : integer := 3082;
        Y3X11           : integer := 3083;
        Y3X12           : integer := 3084;
        Y3X13           : integer := 3085;
        Y3X14           : integer := 3086;
        Y3X15           : integer := 3087;
        Y3X16           : integer := 3088;
        Y3X17           : integer := 3089;
        Y3X18           : integer := 3090;
        Y3X19           : integer := 3091;
        Y3X20           : integer := 3092;
        Y3X21           : integer := 3093;
        Y3X22           : integer := 3094;
        Y3X23           : integer := 3095;
        Y3X24           : integer := 3096;
        Y3X25           : integer := 3097;
        Y3X26           : integer := 3098;
        Y3X27           : integer := 3099;
        Y3X28           : integer := 3100;
        Y4X1            : integer := 4097;
        Y4X2            : integer := 4098;
        Y4X3            : integer := 4099;
        Y4X4            : integer := 4100;
        Y4X5            : integer := 4101;
        Y4X6            : integer := 4102;
        Y4X7            : integer := 4103;
        Y4X8            : integer := 4104;
        Y4X9            : integer := 4105;
        Y4X10           : integer := 4106;
        Y4X11           : integer := 4107;
        Y4X12           : integer := 4108;
        Y4X13           : integer := 4109;
        Y4X14           : integer := 4110;
        Y4X15           : integer := 4111;
        Y4X16           : integer := 4112;
        Y4X17           : integer := 4113;
        Y4X18           : integer := 4114;
        Y4X19           : integer := 4115;
        Y4X20           : integer := 4116;
        Y4X21           : integer := 4117;
        Y4X22           : integer := 4118;
        Y4X23           : integer := 4119;
        Y4X24           : integer := 4120;
        Y4X25           : integer := 4121;
        Y4X26           : integer := 4122;
        Y4X27           : integer := 4123;
        Y4X28           : integer := 4124;
        Y5X1            : integer := 5121;
        Y5X2            : integer := 5122;
        Y5X3            : integer := 5123;
        Y5X4            : integer := 5124;
        Y5X5            : integer := 5125;
        Y5X6            : integer := 5126;
        Y5X7            : integer := 5127;
        Y5X8            : integer := 5128;
        Y5X9            : integer := 5129;
        Y5X10           : integer := 5130;
        Y5X11           : integer := 5131;
        Y5X12           : integer := 5132;
        Y5X13           : integer := 5133;
        Y5X14           : integer := 5134;
        Y5X15           : integer := 5135;
        Y5X16           : integer := 5136;
        Y5X17           : integer := 5137;
        Y5X18           : integer := 5138;
        Y5X19           : integer := 5139;
        Y5X20           : integer := 5140;
        Y5X21           : integer := 5141;
        Y5X22           : integer := 5142;
        Y5X23           : integer := 5143;
        Y5X24           : integer := 5144;
        Y5X25           : integer := 5145;
        Y5X26           : integer := 5146;
        Y5X27           : integer := 5147;
        Y5X28           : integer := 5148;
        Y6X1            : integer := 6145;
        Y6X2            : integer := 6146;
        Y6X3            : integer := 6147;
        Y6X4            : integer := 6148;
        Y6X5            : integer := 6149;
        Y6X6            : integer := 6150;
        Y6X7            : integer := 6151;
        Y6X8            : integer := 6152;
        Y6X9            : integer := 6153;
        Y6X10           : integer := 6154;
        Y6X11           : integer := 6155;
        Y6X12           : integer := 6156;
        Y6X13           : integer := 6157;
        Y6X14           : integer := 6158;
        Y6X15           : integer := 6159;
        Y6X16           : integer := 6160;
        Y6X17           : integer := 6161;
        Y6X18           : integer := 6162;
        Y6X19           : integer := 6163;
        Y6X20           : integer := 6164;
        Y6X21           : integer := 6165;
        Y6X22           : integer := 6166;
        Y6X23           : integer := 6167;
        Y6X24           : integer := 6168;
        Y6X25           : integer := 6169;
        Y6X26           : integer := 6170;
        Y6X27           : integer := 6171;
        Y6X28           : integer := 6172;
        Y7X1            : integer := 7169;
        Y7X2            : integer := 7170;
        Y7X3            : integer := 7171;
        Y7X4            : integer := 7172;
        Y7X5            : integer := 7173;
        Y7X6            : integer := 7174;
        Y7X7            : integer := 7175;
        Y7X8            : integer := 7176;
        Y7X9            : integer := 7177;
        Y7X10           : integer := 7178;
        Y7X11           : integer := 7179;
        Y7X12           : integer := 7180;
        Y7X13           : integer := 7181;
        Y7X14           : integer := 7182;
        Y7X15           : integer := 7183;
        Y7X16           : integer := 7184;
        Y7X17           : integer := 7185;
        Y7X18           : integer := 7186;
        Y7X19           : integer := 7187;
        Y7X20           : integer := 7188;
        Y7X21           : integer := 7189;
        Y7X22           : integer := 7190;
        Y7X23           : integer := 7191;
        Y7X24           : integer := 7192;
        Y7X25           : integer := 7193;
        Y7X26           : integer := 7194;
        Y7X27           : integer := 7195;
        Y7X28           : integer := 7196;
        Y8X1            : integer := 8193;
        Y8X2            : integer := 8194;
        Y8X3            : integer := 8195;
        Y8X4            : integer := 8196;
        Y8X5            : integer := 8197;
        Y8X6            : integer := 8198;
        Y8X7            : integer := 8199;
        Y8X8            : integer := 8200;
        Y8X9            : integer := 8201;
        Y8X10           : integer := 8202;
        Y8X11           : integer := 8203;
        Y8X12           : integer := 8204;
        Y8X13           : integer := 8205;
        Y8X14           : integer := 8206;
        Y8X15           : integer := 8207;
        Y8X16           : integer := 8208;
        Y8X17           : integer := 8209;
        Y8X18           : integer := 8210;
        Y8X19           : integer := 8211;
        Y8X20           : integer := 8212;
        Y8X21           : integer := 8213;
        Y8X22           : integer := 8214;
        Y8X23           : integer := 8215;
        Y8X24           : integer := 8216;
        Y8X25           : integer := 8217;
        Y8X26           : integer := 8218;
        Y8X27           : integer := 8219;
        Y8X28           : integer := 8220;
        Y9X1            : integer := 9217;
        Y9X2            : integer := 9218;
        Y9X3            : integer := 9219;
        Y9X4            : integer := 9220;
        Y9X5            : integer := 9221;
        Y9X6            : integer := 9222;
        Y9X7            : integer := 9223;
        Y9X8            : integer := 9224;
        Y9X9            : integer := 9225;
        Y9X10           : integer := 9226;
        Y9X11           : integer := 9227;
        Y9X12           : integer := 9228;
        Y9X13           : integer := 9229;
        Y9X14           : integer := 9230;
        Y9X15           : integer := 9231;
        Y9X16           : integer := 9232;
        Y9X17           : integer := 9233;
        Y9X18           : integer := 9234;
        Y9X19           : integer := 9235;
        Y9X20           : integer := 9236;
        Y9X21           : integer := 9237;
        Y9X22           : integer := 9238;
        Y9X23           : integer := 9239;
        Y9X24           : integer := 9240;
        Y9X25           : integer := 9241;
        Y9X26           : integer := 9242;
        Y9X27           : integer := 9243;
        Y9X28           : integer := 9244;
        Y10X1           : integer := 10241;
        Y10X2           : integer := 10242;
        Y10X3           : integer := 10243;
        Y10X4           : integer := 10244;
        Y10X5           : integer := 10245;
        Y10X6           : integer := 10246;
        Y10X7           : integer := 10247;
        Y10X8           : integer := 10248;
        Y10X9           : integer := 10249;
        Y10X10          : integer := 10250;
        Y10X11          : integer := 10251;
        Y10X12          : integer := 10252;
        Y10X13          : integer := 10253;
        Y10X14          : integer := 10254;
        Y10X15          : integer := 10255;
        Y10X16          : integer := 10256;
        Y10X17          : integer := 10257;
        Y10X18          : integer := 10258;
        Y10X19          : integer := 10259;
        Y10X20          : integer := 10260;
        Y10X21          : integer := 10261;
        Y10X22          : integer := 10262;
        Y10X23          : integer := 10263;
        Y10X24          : integer := 10264;
        Y10X25          : integer := 10265;
        Y10X26          : integer := 10266;
        Y10X27          : integer := 10267;
        Y10X28          : integer := 10268;
        Y11X1           : integer := 11265;
        Y11X2           : integer := 11266;
        Y11X3           : integer := 11267;
        Y11X4           : integer := 11268;
        Y11X5           : integer := 11269;
        Y11X6           : integer := 11270;
        Y11X7           : integer := 11271;
        Y11X8           : integer := 11272;
        Y11X9           : integer := 11273;
        Y11X10          : integer := 11274;
        Y11X11          : integer := 11275;
        Y11X12          : integer := 11276;
        Y11X13          : integer := 11277;
        Y11X14          : integer := 11278;
        Y11X15          : integer := 11279;
        Y11X16          : integer := 11280;
        Y11X17          : integer := 11281;
        Y11X18          : integer := 11282;
        Y11X19          : integer := 11283;
        Y11X20          : integer := 11284;
        Y11X21          : integer := 11285;
        Y11X22          : integer := 11286;
        Y11X23          : integer := 11287;
        Y11X24          : integer := 11288;
        Y11X25          : integer := 11289;
        Y11X26          : integer := 11290;
        Y11X27          : integer := 11291;
        Y11X28          : integer := 11292;
        Y12X1           : integer := 12289;
        Y12X2           : integer := 12290;
        Y12X3           : integer := 12291;
        Y12X4           : integer := 12292;
        Y12X5           : integer := 12293;
        Y12X6           : integer := 12294;
        Y12X7           : integer := 12295;
        Y12X8           : integer := 12296;
        Y12X9           : integer := 12297;
        Y12X10          : integer := 12298;
        Y12X11          : integer := 12299;
        Y12X12          : integer := 12300;
        Y12X13          : integer := 12301;
        Y12X14          : integer := 12302;
        Y12X15          : integer := 12303;
        Y12X16          : integer := 12304;
        Y12X17          : integer := 12305;
        Y12X18          : integer := 12306;
        Y12X19          : integer := 12307;
        Y12X20          : integer := 12308;
        Y12X21          : integer := 12309;
        Y12X22          : integer := 12310;
        Y12X23          : integer := 12311;
        Y12X24          : integer := 12312;
        Y12X25          : integer := 12313;
        Y12X26          : integer := 12314;
        Y12X27          : integer := 12315;
        Y12X28          : integer := 12316;
        Y13X1           : integer := 13313;
        Y13X2           : integer := 13314;
        Y13X3           : integer := 13315;
        Y13X4           : integer := 13316;
        Y13X5           : integer := 13317;
        Y13X6           : integer := 13318;
        Y13X7           : integer := 13319;
        Y13X8           : integer := 13320;
        Y13X9           : integer := 13321;
        Y13X10          : integer := 13322;
        Y13X11          : integer := 13323;
        Y13X12          : integer := 13324;
        Y13X13          : integer := 13325;
        Y13X14          : integer := 13326;
        Y13X15          : integer := 13327;
        Y13X16          : integer := 13328;
        Y13X17          : integer := 13329;
        Y13X18          : integer := 13330;
        Y13X19          : integer := 13331;
        Y13X20          : integer := 13332;
        Y13X21          : integer := 13333;
        Y13X22          : integer := 13334;
        Y13X23          : integer := 13335;
        Y13X24          : integer := 13336;
        Y13X25          : integer := 13337;
        Y13X26          : integer := 13338;
        Y13X27          : integer := 13339;
        Y13X28          : integer := 13340;
        Y14X1           : integer := 14337;
        Y14X2           : integer := 14338;
        Y14X3           : integer := 14339;
        Y14X4           : integer := 14340;
        Y14X5           : integer := 14341;
        Y14X6           : integer := 14342;
        Y14X7           : integer := 14343;
        Y14X8           : integer := 14344;
        Y14X9           : integer := 14345;
        Y14X10          : integer := 14346;
        Y14X11          : integer := 14347;
        Y14X12          : integer := 14348;
        Y14X13          : integer := 14349;
        Y14X14          : integer := 14350;
        Y14X15          : integer := 14351;
        Y14X16          : integer := 14352;
        Y14X17          : integer := 14353;
        Y14X18          : integer := 14354;
        Y14X19          : integer := 14355;
        Y14X20          : integer := 14356;
        Y14X21          : integer := 14357;
        Y14X22          : integer := 14358;
        Y14X23          : integer := 14359;
        Y14X24          : integer := 14360;
        Y14X25          : integer := 14361;
        Y14X26          : integer := 14362;
        Y14X27          : integer := 14363;
        Y14X28          : integer := 14364;
        Y15X1           : integer := 15361;
        Y15X2           : integer := 15362;
        Y15X3           : integer := 15363;
        Y15X4           : integer := 15364;
        Y15X5           : integer := 15365;
        Y15X6           : integer := 15366;
        Y15X7           : integer := 15367;
        Y15X8           : integer := 15368;
        Y15X9           : integer := 15369;
        Y15X10          : integer := 15370;
        Y15X11          : integer := 15371;
        Y15X12          : integer := 15372;
        Y15X13          : integer := 15373;
        Y15X14          : integer := 15374;
        Y15X15          : integer := 15375;
        Y15X16          : integer := 15376;
        Y15X17          : integer := 15377;
        Y15X18          : integer := 15378;
        Y15X19          : integer := 15379;
        Y15X20          : integer := 15380;
        Y15X21          : integer := 15381;
        Y15X22          : integer := 15382;
        Y15X23          : integer := 15383;
        Y15X24          : integer := 15384;
        Y15X25          : integer := 15385;
        Y15X26          : integer := 15386;
        Y15X27          : integer := 15387;
        Y15X28          : integer := 15388;
        Y16X1           : integer := 16385;
        Y16X2           : integer := 16386;
        Y16X3           : integer := 16387;
        Y16X4           : integer := 16388;
        Y16X5           : integer := 16389;
        Y16X6           : integer := 16390;
        Y16X7           : integer := 16391;
        Y16X8           : integer := 16392;
        Y16X9           : integer := 16393;
        Y16X10          : integer := 16394;
        Y16X11          : integer := 16395;
        Y16X12          : integer := 16396;
        Y16X13          : integer := 16397;
        Y16X14          : integer := 16398;
        Y16X15          : integer := 16399;
        Y16X16          : integer := 16400;
        Y16X17          : integer := 16401;
        Y16X18          : integer := 16402;
        Y16X19          : integer := 16403;
        Y16X20          : integer := 16404;
        Y16X21          : integer := 16405;
        Y16X22          : integer := 16406;
        Y16X23          : integer := 16407;
        Y16X24          : integer := 16408;
        Y16X25          : integer := 16409;
        Y16X26          : integer := 16410;
        Y16X27          : integer := 16411;
        Y16X28          : integer := 16412;
        Y17X1           : integer := 17409;
        Y17X2           : integer := 17410;
        Y17X3           : integer := 17411;
        Y17X4           : integer := 17412;
        Y17X5           : integer := 17413;
        Y17X6           : integer := 17414;
        Y17X7           : integer := 17415;
        Y17X8           : integer := 17416;
        Y17X9           : integer := 17417;
        Y17X10          : integer := 17418;
        Y17X11          : integer := 17419;
        Y17X12          : integer := 17420;
        Y17X13          : integer := 17421;
        Y17X14          : integer := 17422;
        Y17X15          : integer := 17423;
        Y17X16          : integer := 17424;
        Y17X17          : integer := 17425;
        Y17X18          : integer := 17426;
        Y17X19          : integer := 17427;
        Y17X20          : integer := 17428;
        Y17X21          : integer := 17429;
        Y17X22          : integer := 17430;
        Y17X23          : integer := 17431;
        Y17X24          : integer := 17432;
        Y17X25          : integer := 17433;
        Y17X26          : integer := 17434;
        Y17X27          : integer := 17435;
        Y17X28          : integer := 17436;
        Y18X1           : integer := 18433;
        Y18X2           : integer := 18434;
        Y18X3           : integer := 18435;
        Y18X4           : integer := 18436;
        Y18X5           : integer := 18437;
        Y18X6           : integer := 18438;
        Y18X7           : integer := 18439;
        Y18X8           : integer := 18440;
        Y18X9           : integer := 18441;
        Y18X10          : integer := 18442;
        Y18X11          : integer := 18443;
        Y18X12          : integer := 18444;
        Y18X13          : integer := 18445;
        Y18X14          : integer := 18446;
        Y18X15          : integer := 18447;
        Y18X16          : integer := 18448;
        Y18X17          : integer := 18449;
        Y18X18          : integer := 18450;
        Y18X19          : integer := 18451;
        Y18X20          : integer := 18452;
        Y18X21          : integer := 18453;
        Y18X22          : integer := 18454;
        Y18X23          : integer := 18455;
        Y18X24          : integer := 18456;
        Y18X25          : integer := 18457;
        Y18X26          : integer := 18458;
        Y18X27          : integer := 18459;
        Y18X28          : integer := 18460;
        Y19X1           : integer := 19457;
        Y19X2           : integer := 19458;
        Y19X3           : integer := 19459;
        Y19X4           : integer := 19460;
        Y19X5           : integer := 19461;
        Y19X6           : integer := 19462;
        Y19X7           : integer := 19463;
        Y19X8           : integer := 19464;
        Y19X9           : integer := 19465;
        Y19X10          : integer := 19466;
        Y19X11          : integer := 19467;
        Y19X12          : integer := 19468;
        Y19X13          : integer := 19469;
        Y19X14          : integer := 19470;
        Y19X15          : integer := 19471;
        Y19X16          : integer := 19472;
        Y19X17          : integer := 19473;
        Y19X18          : integer := 19474;
        Y19X19          : integer := 19475;
        Y19X20          : integer := 19476;
        Y19X21          : integer := 19477;
        Y19X22          : integer := 19478;
        Y19X23          : integer := 19479;
        Y19X24          : integer := 19480;
        Y19X25          : integer := 19481;
        Y19X26          : integer := 19482;
        Y19X27          : integer := 19483;
        Y19X28          : integer := 19484;
        Y20X1           : integer := 20481;
        Y20X2           : integer := 20482;
        Y20X3           : integer := 20483;
        Y20X4           : integer := 20484;
        Y20X5           : integer := 20485;
        Y20X6           : integer := 20486;
        Y20X7           : integer := 20487;
        Y20X8           : integer := 20488;
        Y20X9           : integer := 20489;
        Y20X10          : integer := 20490;
        Y20X11          : integer := 20491;
        Y20X12          : integer := 20492;
        Y20X13          : integer := 20493;
        Y20X14          : integer := 20494;
        Y20X15          : integer := 20495;
        Y20X16          : integer := 20496;
        Y20X17          : integer := 20497;
        Y20X18          : integer := 20498;
        Y20X19          : integer := 20499;
        Y20X20          : integer := 20500;
        Y20X21          : integer := 20501;
        Y20X22          : integer := 20502;
        Y20X23          : integer := 20503;
        Y20X24          : integer := 20504;
        Y20X25          : integer := 20505;
        Y20X26          : integer := 20506;
        Y20X27          : integer := 20507;
        Y20X28          : integer := 20508;
        Y21X1           : integer := 21505;
        Y21X2           : integer := 21506;
        Y21X3           : integer := 21507;
        Y21X4           : integer := 21508;
        Y21X5           : integer := 21509;
        Y21X6           : integer := 21510;
        Y21X7           : integer := 21511;
        Y21X8           : integer := 21512;
        Y21X9           : integer := 21513;
        Y21X10          : integer := 21514;
        Y21X11          : integer := 21515;
        Y21X12          : integer := 21516;
        Y21X13          : integer := 21517;
        Y21X14          : integer := 21518;
        Y21X15          : integer := 21519;
        Y21X16          : integer := 21520;
        Y21X17          : integer := 21521;
        Y21X18          : integer := 21522;
        Y21X19          : integer := 21523;
        Y21X20          : integer := 21524;
        Y21X21          : integer := 21525;
        Y21X22          : integer := 21526;
        Y21X23          : integer := 21527;
        Y21X24          : integer := 21528;
        Y21X25          : integer := 21529;
        Y21X26          : integer := 21530;
        Y21X27          : integer := 21531;
        Y21X28          : integer := 21532;
        Y22X1           : integer := 22529;
        Y22X2           : integer := 22530;
        Y22X3           : integer := 22531;
        Y22X4           : integer := 22532;
        Y22X5           : integer := 22533;
        Y22X6           : integer := 22534;
        Y22X7           : integer := 22535;
        Y22X8           : integer := 22536;
        Y22X9           : integer := 22537;
        Y22X10          : integer := 22538;
        Y22X11          : integer := 22539;
        Y22X12          : integer := 22540;
        Y22X13          : integer := 22541;
        Y22X14          : integer := 22542;
        Y22X15          : integer := 22543;
        Y22X16          : integer := 22544;
        Y22X17          : integer := 22545;
        Y22X18          : integer := 22546;
        Y22X19          : integer := 22547;
        Y22X20          : integer := 22548;
        Y22X21          : integer := 22549;
        Y22X22          : integer := 22550;
        Y22X23          : integer := 22551;
        Y22X24          : integer := 22552;
        Y22X25          : integer := 22553;
        Y22X26          : integer := 22554;
        Y22X27          : integer := 22555;
        Y22X28          : integer := 22556;
        Y23X1           : integer := 23553;
        Y23X2           : integer := 23554;
        Y23X3           : integer := 23555;
        Y23X4           : integer := 23556;
        Y23X5           : integer := 23557;
        Y23X6           : integer := 23558;
        Y23X7           : integer := 23559;
        Y23X8           : integer := 23560;
        Y23X9           : integer := 23561;
        Y23X10          : integer := 23562;
        Y23X11          : integer := 23563;
        Y23X12          : integer := 23564;
        Y23X13          : integer := 23565;
        Y23X14          : integer := 23566;
        Y23X15          : integer := 23567;
        Y23X16          : integer := 23568;
        Y23X17          : integer := 23569;
        Y23X18          : integer := 23570;
        Y23X19          : integer := 23571;
        Y23X20          : integer := 23572;
        Y23X21          : integer := 23573;
        Y23X22          : integer := 23574;
        Y23X23          : integer := 23575;
        Y23X24          : integer := 23576;
        Y23X25          : integer := 23577;
        Y23X26          : integer := 23578;
        Y23X27          : integer := 23579;
        Y23X28          : integer := 23580;
        Y24X1           : integer := 24577;
        Y24X2           : integer := 24578;
        Y24X3           : integer := 24579;
        Y24X4           : integer := 24580;
        Y24X5           : integer := 24581;
        Y24X6           : integer := 24582;
        Y24X7           : integer := 24583;
        Y24X8           : integer := 24584;
        Y24X9           : integer := 24585;
        Y24X10          : integer := 24586;
        Y24X11          : integer := 24587;
        Y24X12          : integer := 24588;
        Y24X13          : integer := 24589;
        Y24X14          : integer := 24590;
        Y24X15          : integer := 24591;
        Y24X16          : integer := 24592;
        Y24X17          : integer := 24593;
        Y24X18          : integer := 24594;
        Y24X19          : integer := 24595;
        Y24X20          : integer := 24596;
        Y24X21          : integer := 24597;
        Y24X22          : integer := 24598;
        Y24X23          : integer := 24599;
        Y24X24          : integer := 24600;
        Y24X25          : integer := 24601;
        Y24X26          : integer := 24602;
        Y24X27          : integer := 24603;
        Y24X28          : integer := 24604;
        Y25X1           : integer := 25601;
        Y25X2           : integer := 25602;
        Y25X3           : integer := 25603;
        Y25X4           : integer := 25604;
        Y25X5           : integer := 25605;
        Y25X6           : integer := 25606;
        Y25X7           : integer := 25607;
        Y25X8           : integer := 25608;
        Y25X9           : integer := 25609;
        Y25X10          : integer := 25610;
        Y25X11          : integer := 25611;
        Y25X12          : integer := 25612;
        Y25X13          : integer := 25613;
        Y25X14          : integer := 25614;
        Y25X15          : integer := 25615;
        Y25X16          : integer := 25616;
        Y25X17          : integer := 25617;
        Y25X18          : integer := 25618;
        Y25X19          : integer := 25619;
        Y25X20          : integer := 25620;
        Y25X21          : integer := 25621;
        Y25X22          : integer := 25622;
        Y25X23          : integer := 25623;
        Y25X24          : integer := 25624;
        Y25X25          : integer := 25625;
        Y25X26          : integer := 25626;
        Y25X27          : integer := 25627;
        Y25X28          : integer := 25628;
        Y26X1           : integer := 26625;
        Y26X2           : integer := 26626;
        Y26X3           : integer := 26627;
        Y26X4           : integer := 26628;
        Y26X5           : integer := 26629;
        Y26X6           : integer := 26630;
        Y26X7           : integer := 26631;
        Y26X8           : integer := 26632;
        Y26X9           : integer := 26633;
        Y26X10          : integer := 26634;
        Y26X11          : integer := 26635;
        Y26X12          : integer := 26636;
        Y26X13          : integer := 26637;
        Y26X14          : integer := 26638;
        Y26X15          : integer := 26639;
        Y26X16          : integer := 26640;
        Y26X17          : integer := 26641;
        Y26X18          : integer := 26642;
        Y26X19          : integer := 26643;
        Y26X20          : integer := 26644;
        Y26X21          : integer := 26645;
        Y26X22          : integer := 26646;
        Y26X23          : integer := 26647;
        Y26X24          : integer := 26648;
        Y26X25          : integer := 26649;
        Y26X26          : integer := 26650;
        Y26X27          : integer := 26651;
        Y26X28          : integer := 26652;
        Y27X1           : integer := 27649;
        Y27X2           : integer := 27650;
        Y27X3           : integer := 27651;
        Y27X4           : integer := 27652;
        Y27X5           : integer := 27653;
        Y27X6           : integer := 27654;
        Y27X7           : integer := 27655;
        Y27X8           : integer := 27656;
        Y27X9           : integer := 27657;
        Y27X10          : integer := 27658;
        Y27X11          : integer := 27659;
        Y27X12          : integer := 27660;
        Y27X13          : integer := 27661;
        Y27X14          : integer := 27662;
        Y27X15          : integer := 27663;
        Y27X16          : integer := 27664;
        Y27X17          : integer := 27665;
        Y27X18          : integer := 27666;
        Y27X19          : integer := 27667;
        Y27X20          : integer := 27668;
        Y27X21          : integer := 27669;
        Y27X22          : integer := 27670;
        Y27X23          : integer := 27671;
        Y27X24          : integer := 27672;
        Y27X25          : integer := 27673;
        Y27X26          : integer := 27674;
        Y27X27          : integer := 27675;
        Y27X28          : integer := 27676;
        Y28X1           : integer := 28673;
        Y28X2           : integer := 28674;
        Y28X3           : integer := 28675;
        Y28X4           : integer := 28676;
        Y28X5           : integer := 28677;
        Y28X6           : integer := 28678;
        Y28X7           : integer := 28679;
        Y28X8           : integer := 28680;
        Y28X9           : integer := 28681;
        Y28X10          : integer := 28682;
        Y28X11          : integer := 28683;
        Y28X12          : integer := 28684;
        Y28X13          : integer := 28685;
        Y28X14          : integer := 28686;
        Y28X15          : integer := 28687;
        Y28X16          : integer := 28688;
        Y28X17          : integer := 28689;
        Y28X18          : integer := 28690;
        Y28X19          : integer := 28691;
        Y28X20          : integer := 28692;
        Y28X21          : integer := 28693;
        Y28X22          : integer := 28694;
        Y28X23          : integer := 28695;
        Y28X24          : integer := 28696;
        Y28X25          : integer := 28697;
        Y28X26          : integer := 28698;
        Y28X27          : integer := 28699;
        Y28X28          : integer := 28700;
        Y29X1           : integer := 29697;
        Y29X2           : integer := 29698;
        Y29X3           : integer := 29699;
        Y29X4           : integer := 29700;
        Y29X5           : integer := 29701;
        Y29X6           : integer := 29702;
        Y29X7           : integer := 29703;
        Y29X8           : integer := 29704;
        Y29X9           : integer := 29705;
        Y29X10          : integer := 29706;
        Y29X11          : integer := 29707;
        Y29X12          : integer := 29708;
        Y29X13          : integer := 29709;
        Y29X14          : integer := 29710;
        Y29X15          : integer := 29711;
        Y29X16          : integer := 29712;
        Y29X17          : integer := 29713;
        Y29X18          : integer := 29714;
        Y29X19          : integer := 29715;
        Y29X20          : integer := 29716;
        Y29X21          : integer := 29717;
        Y29X22          : integer := 29718;
        Y29X23          : integer := 29719;
        Y29X24          : integer := 29720;
        Y29X25          : integer := 29721;
        Y29X26          : integer := 29722;
        Y29X27          : integer := 29723;
        Y29X28          : integer := 29724;
        Y30X1           : integer := 30721;
        Y30X2           : integer := 30722;
        Y30X3           : integer := 30723;
        Y30X4           : integer := 30724;
        Y30X5           : integer := 30725;
        Y30X6           : integer := 30726;
        Y30X7           : integer := 30727;
        Y30X8           : integer := 30728;
        Y30X9           : integer := 30729;
        Y30X10          : integer := 30730;
        Y30X11          : integer := 30731;
        Y30X12          : integer := 30732;
        Y30X13          : integer := 30733;
        Y30X14          : integer := 30734;
        Y30X15          : integer := 30735;
        Y30X16          : integer := 30736;
        Y30X17          : integer := 30737;
        Y30X18          : integer := 30738;
        Y30X19          : integer := 30739;
        Y30X20          : integer := 30740;
        Y30X21          : integer := 30741;
        Y30X22          : integer := 30742;
        Y30X23          : integer := 30743;
        Y30X24          : integer := 30744;
        Y30X25          : integer := 30745;
        Y30X26          : integer := 30746;
        Y30X27          : integer := 30747;
        Y30X28          : integer := 30748;
        Y31X1           : integer := 31745;
        Y31X2           : integer := 31746;
        Y31X3           : integer := 31747;
        Y31X4           : integer := 31748;
        Y31X5           : integer := 31749;
        Y31X6           : integer := 31750;
        Y31X7           : integer := 31751;
        Y31X8           : integer := 31752;
        Y31X9           : integer := 31753;
        Y31X10          : integer := 31754;
        Y31X11          : integer := 31755;
        Y31X12          : integer := 31756;
        Y31X13          : integer := 31757;
        Y31X14          : integer := 31758;
        Y31X15          : integer := 31759;
        Y31X16          : integer := 31760;
        Y31X17          : integer := 31761;
        Y31X18          : integer := 31762;
        Y31X19          : integer := 31763;
        Y31X20          : integer := 31764;
        Y31X21          : integer := 31765;
        Y31X22          : integer := 31766;
        Y31X23          : integer := 31767;
        Y31X24          : integer := 31768;
        Y31X25          : integer := 31769;
        Y31X26          : integer := 31770;
        Y31X27          : integer := 31771;
        Y31X28          : integer := 31772;
        Y32X1           : integer := 32769;
        Y32X2           : integer := 32770;
        Y32X3           : integer := 32771;
        Y32X4           : integer := 32772;
        Y32X5           : integer := 32773;
        Y32X6           : integer := 32774;
        Y32X7           : integer := 32775;
        Y32X8           : integer := 32776;
        Y32X9           : integer := 32777;
        Y32X10          : integer := 32778;
        Y32X11          : integer := 32779;
        Y32X12          : integer := 32780;
        Y32X13          : integer := 32781;
        Y32X14          : integer := 32782;
        Y32X15          : integer := 32783;
        Y32X16          : integer := 32784;
        Y32X17          : integer := 32785;
        Y32X18          : integer := 32786;
        Y32X19          : integer := 32787;
        Y32X20          : integer := 32788;
        Y32X21          : integer := 32789;
        Y32X22          : integer := 32790;
        Y32X23          : integer := 32791;
        Y32X24          : integer := 32792;
        Y32X25          : integer := 32793;
        Y32X26          : integer := 32794;
        Y32X27          : integer := 32795;
        Y32X28          : integer := 32796;
        Y33X1           : integer := 33793;
        Y33X2           : integer := 33794;
        Y33X3           : integer := 33795;
        Y33X4           : integer := 33796;
        Y33X5           : integer := 33797;
        Y33X6           : integer := 33798;
        Y33X7           : integer := 33799;
        Y33X8           : integer := 33800;
        Y33X9           : integer := 33801;
        Y33X10          : integer := 33802;
        Y33X11          : integer := 33803;
        Y33X12          : integer := 33804;
        Y33X13          : integer := 33805;
        Y33X14          : integer := 33806;
        Y33X15          : integer := 33807;
        Y33X16          : integer := 33808;
        Y33X17          : integer := 33809;
        Y33X18          : integer := 33810;
        Y33X19          : integer := 33811;
        Y33X20          : integer := 33812;
        Y33X21          : integer := 33813;
        Y33X22          : integer := 33814;
        Y33X23          : integer := 33815;
        Y33X24          : integer := 33816;
        Y33X25          : integer := 33817;
        Y33X26          : integer := 33818;
        Y33X27          : integer := 33819;
        Y33X28          : integer := 33820;
        Y34X1           : integer := 34817;
        Y34X2           : integer := 34818;
        Y34X3           : integer := 34819;
        Y34X4           : integer := 34820;
        Y34X5           : integer := 34821;
        Y34X6           : integer := 34822;
        Y34X7           : integer := 34823;
        Y34X8           : integer := 34824;
        Y34X9           : integer := 34825;
        Y34X10          : integer := 34826;
        Y34X11          : integer := 34827;
        Y34X12          : integer := 34828;
        Y34X13          : integer := 34829;
        Y34X14          : integer := 34830;
        Y34X15          : integer := 34831;
        Y34X16          : integer := 34832;
        Y34X17          : integer := 34833;
        Y34X18          : integer := 34834;
        Y34X19          : integer := 34835;
        Y34X20          : integer := 34836;
        Y34X21          : integer := 34837;
        Y34X22          : integer := 34838;
        Y34X23          : integer := 34839;
        Y34X24          : integer := 34840;
        Y34X25          : integer := 34841;
        Y34X26          : integer := 34842;
        Y34X27          : integer := 34843;
        Y34X28          : integer := 34844;
        Y35X1           : integer := 35841;
        Y35X2           : integer := 35842;
        Y35X3           : integer := 35843;
        Y35X4           : integer := 35844;
        Y35X5           : integer := 35845;
        Y35X6           : integer := 35846;
        Y35X7           : integer := 35847;
        Y35X8           : integer := 35848;
        Y35X9           : integer := 35849;
        Y35X10          : integer := 35850;
        Y35X11          : integer := 35851;
        Y35X12          : integer := 35852;
        Y35X13          : integer := 35853;
        Y35X14          : integer := 35854;
        Y35X15          : integer := 35855;
        Y35X16          : integer := 35856;
        Y35X17          : integer := 35857;
        Y35X18          : integer := 35858;
        Y35X19          : integer := 35859;
        Y35X20          : integer := 35860;
        Y35X21          : integer := 35861;
        Y35X22          : integer := 35862;
        Y35X23          : integer := 35863;
        Y35X24          : integer := 35864;
        Y35X25          : integer := 35865;
        Y35X26          : integer := 35866;
        Y35X27          : integer := 35867;
        Y35X28          : integer := 35868;
        YY0XX0          : integer := 3840;
        YY0XX1          : integer := 819;
        YY0XX2          : integer := 1621;
        YY0XX3          : integer := 1637;
        YY0XX4          : integer := 1910;
        YY0XX5          : integer := 3840;
        YY0XX6          : integer := 3840;
        YY0XX7          : integer := 3840;
        YY0XX8          : integer := 3840;
        YY0XX9          : integer := 3840;
        YY0XX10         : integer := 3840;
        YY0XX11         : integer := 3840;
        YY0XX12         : integer := 3840;
        YY0XX13         : integer := 3840;
        YY0XX14         : integer := 3840;
        YY0XX15         : integer := 3840;
        YY0XX16         : integer := 3840;
        YY0XX17         : integer := 3840;
        YY0XX18         : integer := 3840;
        YY0XX19         : integer := 3840;
        YY0XX20         : integer := 3840;
        YY0XX21         : integer := 3840;
        YY0XX22         : integer := 3840;
        YY0XX23         : integer := 3840;
        YY0XX24         : integer := 3840;
        YY0XX25         : integer := 3840;
        YY0XX26         : integer := 3840;
        YY0XX27         : integer := 3840;
        YY0XX28         : integer := 3840;
        YY1XX1          : integer := 2184;
        YY1XX2          : integer := 3276;
        YY1XX3          : integer := 3532;
        YY1XX4          : integer := 3549;
        YY1XX5          : integer := 3002;
        YY1XX6          : integer := 2183;
        YY1XX7          : integer := 3840;
        YY1XX8          : integer := 3840;
        YY1XX9          : integer := 3840;
        YY1XX10         : integer := 3840;
        YY1XX11         : integer := 3840;
        YY1XX12         : integer := 3840;
        YY1XX13         : integer := 3840;
        YY1XX14         : integer := 3840;
        YY1XX15         : integer := 3840;
        YY1XX16         : integer := 3840;
        YY1XX17         : integer := 3840;
        YY1XX18         : integer := 3840;
        YY1XX19         : integer := 3840;
        YY1XX20         : integer := 3840;
        YY1XX21         : integer := 3840;
        YY1XX22         : integer := 3840;
        YY1XX23         : integer := 3840;
        YY1XX24         : integer := 3840;
        YY1XX25         : integer := 3840;
        YY1XX26         : integer := 3840;
        YY1XX27         : integer := 3840;
        YY1XX28         : integer := 3840;
        YY2XX1          : integer := 3003;
        YY2XX2          : integer := 4095;
        YY2XX3          : integer := 4095;
        YY2XX4          : integer := 4095;
        YY2XX5          : integer := 4095;
        YY2XX6          : integer := 3805;
        YY2XX7          : integer := 2713;
        YY2XX8          : integer := 3840;
        YY2XX9          : integer := 3840;
        YY2XX10         : integer := 3840;
        YY2XX11         : integer := 3840;
        YY2XX12         : integer := 3840;
        YY2XX13         : integer := 3840;
        YY2XX14         : integer := 3840;
        YY2XX15         : integer := 3840;
        YY2XX16         : integer := 3840;
        YY2XX17         : integer := 3840;
        YY2XX18         : integer := 3840;
        YY2XX19         : integer := 3840;
        YY2XX20         : integer := 3840;
        YY2XX21         : integer := 3840;
        YY2XX22         : integer := 3840;
        YY2XX23         : integer := 3840;
        YY2XX24         : integer := 3840;
        YY2XX25         : integer := 3840;
        YY2XX26         : integer := 3840;
        YY2XX27         : integer := 3840;
        YY2XX28         : integer := 3840;
        YY3XX1          : integer := 3003;
        YY3XX2          : integer := 4095;
        YY3XX3          : integer := 4095;
        YY3XX4          : integer := 4095;
        YY3XX5          : integer := 4095;
        YY3XX6          : integer := 4095;
        YY3XX7          : integer := 4079;
        YY3XX8          : integer := 3259;
        YY3XX9          : integer := 3840;
        YY3XX10         : integer := 3840;
        YY3XX11         : integer := 3840;
        YY3XX12         : integer := 3840;
        YY3XX13         : integer := 3840;
        YY3XX14         : integer := 3840;
        YY3XX15         : integer := 3840;
        YY3XX16         : integer := 3840;
        YY3XX17         : integer := 3840;
        YY3XX18         : integer := 3840;
        YY3XX19         : integer := 3840;
        YY3XX20         : integer := 3840;
        YY3XX21         : integer := 3840;
        YY3XX22         : integer := 3840;
        YY3XX23         : integer := 3840;
        YY3XX24         : integer := 3840;
        YY3XX25         : integer := 3840;
        YY3XX26         : integer := 3840;
        YY3XX27         : integer := 3840;
        YY3XX28         : integer := 3840;
        YY4XX1          : integer := 2730;
        YY4XX2          : integer := 3550;
        YY4XX3          : integer := 4095;
        YY4XX4          : integer := 4095;
        YY4XX5          : integer := 4095;
        YY4XX6          : integer := 4095;
        YY4XX7          : integer := 4095;
        YY4XX8          : integer := 4095;
        YY4XX9          : integer := 3531;
        YY4XX10         : integer := 3840;
        YY4XX11         : integer := 3840;
        YY4XX12         : integer := 3840;
        YY4XX13         : integer := 3840;
        YY4XX14         : integer := 3840;
        YY4XX15         : integer := 3840;
        YY4XX16         : integer := 3840;
        YY4XX17         : integer := 3840;
        YY4XX18         : integer := 3840;
        YY4XX19         : integer := 3840;
        YY4XX20         : integer := 3840;
        YY4XX21         : integer := 3840;
        YY4XX22         : integer := 3840;
        YY4XX23         : integer := 3840;
        YY4XX24         : integer := 3840;
        YY4XX25         : integer := 3840;
        YY4XX26         : integer := 3840;
        YY4XX27         : integer := 3840;
        YY4XX28         : integer := 3840;
        YY5XX1          : integer := 1927;
        YY5XX2          : integer := 3003;
        YY5XX3          : integer := 3822;
        YY5XX4          : integer := 4095;
        YY5XX5          : integer := 4095;
        YY5XX6          : integer := 4095;
        YY5XX7          : integer := 4095;
        YY5XX8          : integer := 4095;
        YY5XX9          : integer := 4095;
        YY5XX10         : integer := 3532;
        YY5XX11         : integer := 3840;
        YY5XX12         : integer := 3840;
        YY5XX13         : integer := 3840;
        YY5XX14         : integer := 3840;
        YY5XX15         : integer := 3840;
        YY5XX16         : integer := 3840;
        YY5XX17         : integer := 3840;
        YY5XX18         : integer := 3840;
        YY5XX19         : integer := 3840;
        YY5XX20         : integer := 3840;
        YY5XX21         : integer := 3840;
        YY5XX22         : integer := 3840;
        YY5XX23         : integer := 3840;
        YY5XX24         : integer := 3840;
        YY5XX25         : integer := 3840;
        YY5XX26         : integer := 3840;
        YY5XX27         : integer := 3840;
        YY5XX28         : integer := 3840;
        YY6XX1          : integer := 1365;
        YY6XX2          : integer := 2201;
        YY6XX3          : integer := 3276;
        YY6XX4          : integer := 4095;
        YY6XX5          : integer := 4095;
        YY6XX6          : integer := 4095;
        YY6XX7          : integer := 4095;
        YY6XX8          : integer := 4095;
        YY6XX9          : integer := 4095;
        YY6XX10         : integer := 4079;
        YY6XX11         : integer := 3533;
        YY6XX12         : integer := 2730;
        YY6XX13         : integer := 3840;
        YY6XX14         : integer := 3840;
        YY6XX15         : integer := 3840;
        YY6XX16         : integer := 3840;
        YY6XX17         : integer := 3840;
        YY6XX18         : integer := 3840;
        YY6XX19         : integer := 1075;
        YY6XX20         : integer := 1075;
        YY6XX21         : integer := 818;
        YY6XX22         : integer := 3840;
        YY6XX23         : integer := 3840;
        YY6XX24         : integer := 3840;
        YY6XX25         : integer := 3840;
        YY6XX26         : integer := 3840;
        YY6XX27         : integer := 3840;
        YY6XX28         : integer := 3840;
        YY7XX1          : integer := 3840;
        YY7XX2          : integer := 1365;
        YY7XX3          : integer := 2185;
        YY7XX4          : integer := 3276;
        YY7XX5          : integer := 3822;
        YY7XX6          : integer := 4095;
        YY7XX7          : integer := 4095;
        YY7XX8          : integer := 4095;
        YY7XX9          : integer := 4095;
        YY7XX10         : integer := 4095;
        YY7XX11         : integer := 4095;
        YY7XX12         : integer := 4078;
        YY7XX13         : integer := 3003;
        YY7XX14         : integer := 3840;
        YY7XX15         : integer := 3840;
        YY7XX16         : integer := 3840;
        YY7XX17         : integer := 3840;
        YY7XX18         : integer := 1894;
        YY7XX19         : integer := 2456;
        YY7XX20         : integer := 2713;
        YY7XX21         : integer := 1911;
        YY7XX22         : integer := 1091;
        YY7XX23         : integer := 3840;
        YY7XX24         : integer := 3840;
        YY7XX25         : integer := 3840;
        YY7XX26         : integer := 3840;
        YY7XX27         : integer := 3840;
        YY7XX28         : integer := 3840;
        YY8XX1          : integer := 3840;
        YY8XX2          : integer := 3840;
        YY8XX3          : integer := 1092;
        YY8XX4          : integer := 2168;
        YY8XX5          : integer := 2987;
        YY8XX6          : integer := 3822;
        YY8XX7          : integer := 4095;
        YY8XX8          : integer := 4095;
        YY8XX9          : integer := 4095;
        YY8XX10         : integer := 4095;
        YY8XX11         : integer := 4095;
        YY8XX12         : integer := 4095;
        YY8XX13         : integer := 3822;
        YY8XX14         : integer := 3259;
        YY8XX15         : integer := 2440;
        YY8XX16         : integer := 1911;
        YY8XX17         : integer := 1894;
        YY8XX18         : integer := 2440;
        YY8XX19         : integer := 3532;
        YY8XX20         : integer := 4078;
        YY8XX21         : integer := 3275;
        YY8XX22         : integer := 2167;
        YY8XX23         : integer := 2439;
        YY8XX24         : integer := 3840;
        YY8XX25         : integer := 3840;
        YY8XX26         : integer := 3840;
        YY8XX27         : integer := 3840;
        YY8XX28         : integer := 3840;
        YY9XX1          : integer := 3840;
        YY9XX2          : integer := 3840;
        YY9XX3          : integer := 3840;
        YY9XX4          : integer := 1076;
        YY9XX5          : integer := 1895;
        YY9XX6          : integer := 2987;
        YY9XX7          : integer := 3822;
        YY9XX8          : integer := 4095;
        YY9XX9          : integer := 4095;
        YY9XX10         : integer := 4095;
        YY9XX11         : integer := 4095;
        YY9XX12         : integer := 4095;
        YY9XX13         : integer := 4095;
        YY9XX14         : integer := 4095;
        YY9XX15         : integer := 3549;
        YY9XX16         : integer := 3259;
        YY9XX17         : integer := 2730;
        YY9XX18         : integer := 2986;
        YY9XX19         : integer := 3805;
        YY9XX20         : integer := 4095;
        YY9XX21         : integer := 4078;
        YY9XX22         : integer := 3275;
        YY9XX23         : integer := 2439;
        YY9XX24         : integer := 2166;
        YY9XX25         : integer := 3840;
        YY9XX26         : integer := 3840;
        YY9XX27         : integer := 3840;
        YY9XX28         : integer := 3840;
        YY10XX1         : integer := 3840;
        YY10XX2         : integer := 3840;
        YY10XX3         : integer := 3840;
        YY10XX4         : integer := 3840;
        YY10XX5         : integer := 1349;
        YY10XX6         : integer := 2168;
        YY10XX7         : integer := 3003;
        YY10XX8         : integer := 3549;
        YY10XX9         : integer := 4095;
        YY10XX10        : integer := 4095;
        YY10XX11        : integer := 4095;
        YY10XX12        : integer := 4095;
        YY10XX13        : integer := 4095;
        YY10XX14        : integer := 4095;
        YY10XX15        : integer := 4095;
        YY10XX16        : integer := 4095;
        YY10XX17        : integer := 3822;
        YY10XX18        : integer := 3549;
        YY10XX19        : integer := 3805;
        YY10XX20        : integer := 4095;
        YY10XX21        : integer := 4095;
        YY10XX22        : integer := 4095;
        YY10XX23        : integer := 3258;
        YY10XX24        : integer := 2439;
        YY10XX25        : integer := 3840;
        YY10XX26        : integer := 3840;
        YY10XX27        : integer := 3840;
        YY10XX28        : integer := 3840;
        YY11XX1         : integer := 3840;
        YY11XX2         : integer := 3840;
        YY11XX3         : integer := 3840;
        YY11XX4         : integer := 1076;
        YY11XX5         : integer := 1622;
        YY11XX6         : integer := 2457;
        YY11XX7         : integer := 3260;
        YY11XX8         : integer := 3549;
        YY11XX9         : integer := 4095;
        YY11XX10        : integer := 4095;
        YY11XX11        : integer := 4095;
        YY11XX12        : integer := 4095;
        YY11XX13        : integer := 4095;
        YY11XX14        : integer := 4095;
        YY11XX15        : integer := 4095;
        YY11XX16        : integer := 4095;
        YY11XX17        : integer := 4095;
        YY11XX18        : integer := 3822;
        YY11XX19        : integer := 3806;
        YY11XX20        : integer := 3822;
        YY11XX21        : integer := 4095;
        YY11XX22        : integer := 4095;
        YY11XX23        : integer := 4094;
        YY11XX24        : integer := 3531;
        YY11XX25        : integer := 1893;
        YY11XX26        : integer := 3840;
        YY11XX27        : integer := 3840;
        YY11XX28        : integer := 3840;
        YY12XX1         : integer := 3840;
        YY12XX2         : integer := 3840;
        YY12XX3         : integer := 803;
        YY12XX4         : integer := 1365;
        YY12XX5         : integer := 2184;
        YY12XX6         : integer := 3276;
        YY12XX7         : integer := 4079;
        YY12XX8         : integer := 4079;
        YY12XX9         : integer := 4095;
        YY12XX10        : integer := 4095;
        YY12XX11        : integer := 4095;
        YY12XX12        : integer := 4095;
        YY12XX13        : integer := 4095;
        YY12XX14        : integer := 4095;
        YY12XX15        : integer := 4095;
        YY12XX16        : integer := 4095;
        YY12XX17        : integer := 4095;
        YY12XX18        : integer := 4095;
        YY12XX19        : integer := 4095;
        YY12XX20        : integer := 4095;
        YY12XX21        : integer := 4095;
        YY12XX22        : integer := 4095;
        YY12XX23        : integer := 4095;
        YY12XX24        : integer := 4094;
        YY12XX25        : integer := 2729;
        YY12XX26        : integer := 3840;
        YY12XX27        : integer := 3840;
        YY12XX28        : integer := 3840;
        YY13XX1         : integer := 3840;
        YY13XX2         : integer := 3840;
        YY13XX3         : integer := 1638;
        YY13XX4         : integer := 2457;
        YY13XX5         : integer := 3276;
        YY13XX6         : integer := 3822;
        YY13XX7         : integer := 4095;
        YY13XX8         : integer := 4095;
        YY13XX9         : integer := 4095;
        YY13XX10        : integer := 4095;
        YY13XX11        : integer := 4095;
        YY13XX12        : integer := 4095;
        YY13XX13        : integer := 4095;
        YY13XX14        : integer := 4095;
        YY13XX15        : integer := 4095;
        YY13XX16        : integer := 4095;
        YY13XX17        : integer := 4095;
        YY13XX18        : integer := 4095;
        YY13XX19        : integer := 4095;
        YY13XX20        : integer := 4095;
        YY13XX21        : integer := 4095;
        YY13XX22        : integer := 4095;
        YY13XX23        : integer := 4095;
        YY13XX24        : integer := 4078;
        YY13XX25        : integer := 2985;
        YY13XX26        : integer := 3840;
        YY13XX27        : integer := 3840;
        YY13XX28        : integer := 3840;
        YY14XX1         : integer := 3840;
        YY14XX2         : integer := 1365;
        YY14XX3         : integer := 2184;
        YY14XX4         : integer := 3276;
        YY14XX5         : integer := 3822;
        YY14XX6         : integer := 4095;
        YY14XX7         : integer := 4095;
        YY14XX8         : integer := 4095;
        YY14XX9         : integer := 4095;
        YY14XX10        : integer := 4095;
        YY14XX11        : integer := 4095;
        YY14XX12        : integer := 4095;
        YY14XX13        : integer := 4095;
        YY14XX14        : integer := 4095;
        YY14XX15        : integer := 4095;
        YY14XX16        : integer := 4095;
        YY14XX17        : integer := 4095;
        YY14XX18        : integer := 4095;
        YY14XX19        : integer := 4095;
        YY14XX20        : integer := 4095;
        YY14XX21        : integer := 4095;
        YY14XX22        : integer := 4095;
        YY14XX23        : integer := 4095;
        YY14XX24        : integer := 4094;
        YY14XX25        : integer := 2986;
        YY14XX26        : integer := 3840;
        YY14XX27        : integer := 3840;
        YY14XX28        : integer := 3840;
        YY15XX1         : integer := 3840;
        YY15XX2         : integer := 1637;
        YY15XX3         : integer := 2473;
        YY15XX4         : integer := 3565;
        YY15XX5         : integer := 4095;
        YY15XX6         : integer := 4095;
        YY15XX7         : integer := 4095;
        YY15XX8         : integer := 4095;
        YY15XX9         : integer := 4095;
        YY15XX10        : integer := 4095;
        YY15XX11        : integer := 4095;
        YY15XX12        : integer := 4095;
        YY15XX13        : integer := 4095;
        YY15XX14        : integer := 4095;
        YY15XX15        : integer := 4095;
        YY15XX16        : integer := 4095;
        YY15XX17        : integer := 4095;
        YY15XX18        : integer := 4095;
        YY15XX19        : integer := 4095;
        YY15XX20        : integer := 4095;
        YY15XX21        : integer := 4095;
        YY15XX22        : integer := 4095;
        YY15XX23        : integer := 4095;
        YY15XX24        : integer := 4094;
        YY15XX25        : integer := 2713;
        YY15XX26        : integer := 3840;
        YY15XX27        : integer := 3840;
        YY15XX28        : integer := 3840;
        YY16XX1         : integer := 3840;
        YY16XX2         : integer := 1364;
        YY16XX3         : integer := 2456;
        YY16XX4         : integer := 3565;
        YY16XX5         : integer := 3839;
        YY16XX6         : integer := 4095;
        YY16XX7         : integer := 4095;
        YY16XX8         : integer := 4095;
        YY16XX9         : integer := 4095;
        YY16XX10        : integer := 4095;
        YY16XX11        : integer := 4095;
        YY16XX12        : integer := 4095;
        YY16XX13        : integer := 4095;
        YY16XX14        : integer := 4095;
        YY16XX15        : integer := 4095;
        YY16XX16        : integer := 4095;
        YY16XX17        : integer := 4095;
        YY16XX18        : integer := 4095;
        YY16XX19        : integer := 4095;
        YY16XX20        : integer := 4095;
        YY16XX21        : integer := 4095;
        YY16XX22        : integer := 4095;
        YY16XX23        : integer := 4095;
        YY16XX24        : integer := 3822;
        YY16XX25        : integer := 2456;
        YY16XX26        : integer := 3840;
        YY16XX27        : integer := 3840;
        YY16XX28        : integer := 3840;
        YY17XX1         : integer := 3840;
        YY17XX2         : integer := 1075;
        YY17XX3         : integer := 2183;
        YY17XX4         : integer := 3549;
        YY17XX5         : integer := 3839;
        YY17XX6         : integer := 4095;
        YY17XX7         : integer := 4095;
        YY17XX8         : integer := 4095;
        YY17XX9         : integer := 4095;
        YY17XX10        : integer := 4095;
        YY17XX11        : integer := 4095;
        YY17XX12        : integer := 4095;
        YY17XX13        : integer := 4095;
        YY17XX14        : integer := 4095;
        YY17XX15        : integer := 4095;
        YY17XX16        : integer := 4095;
        YY17XX17        : integer := 4095;
        YY17XX18        : integer := 4095;
        YY17XX19        : integer := 4095;
        YY17XX20        : integer := 4095;
        YY17XX21        : integer := 4095;
        YY17XX22        : integer := 4095;
        YY17XX23        : integer := 4095;
        YY17XX24        : integer := 3822;
        YY17XX25        : integer := 2184;
        YY17XX26        : integer := 3840;
        YY17XX27        : integer := 3840;
        YY17XX28        : integer := 3840;
        YY18XX1         : integer := 3840;
        YY18XX2         : integer := 1364;
        YY18XX3         : integer := 2456;
        YY18XX4         : integer := 3549;
        YY18XX5         : integer := 3822;
        YY18XX6         : integer := 4095;
        YY18XX7         : integer := 4095;
        YY18XX8         : integer := 4095;
        YY18XX9         : integer := 4095;
        YY18XX10        : integer := 4095;
        YY18XX11        : integer := 4095;
        YY18XX12        : integer := 4095;
        YY18XX13        : integer := 4095;
        YY18XX14        : integer := 4095;
        YY18XX15        : integer := 4095;
        YY18XX16        : integer := 4095;
        YY18XX17        : integer := 4095;
        YY18XX18        : integer := 4095;
        YY18XX19        : integer := 4095;
        YY18XX20        : integer := 4095;
        YY18XX21        : integer := 4095;
        YY18XX22        : integer := 4095;
        YY18XX23        : integer := 4095;
        YY18XX24        : integer := 3822;
        YY18XX25        : integer := 2184;
        YY18XX26        : integer := 3840;
        YY18XX27        : integer := 3840;
        YY18XX28        : integer := 3840;
        YY19XX1         : integer := 1619;
        YY19XX2         : integer := 2439;
        YY19XX3         : integer := 3003;
        YY19XX4         : integer := 3805;
        YY19XX5         : integer := 3822;
        YY19XX6         : integer := 4095;
        YY19XX7         : integer := 4095;
        YY19XX8         : integer := 4095;
        YY19XX9         : integer := 4095;
        YY19XX10        : integer := 4095;
        YY19XX11        : integer := 4095;
        YY19XX12        : integer := 4095;
        YY19XX13        : integer := 4095;
        YY19XX14        : integer := 4095;
        YY19XX15        : integer := 4095;
        YY19XX16        : integer := 4095;
        YY19XX17        : integer := 4095;
        YY19XX18        : integer := 4095;
        YY19XX19        : integer := 4095;
        YY19XX20        : integer := 4095;
        YY19XX21        : integer := 4095;
        YY19XX22        : integer := 4095;
        YY19XX23        : integer := 4095;
        YY19XX24        : integer := 3565;
        YY19XX25        : integer := 2183;
        YY19XX26        : integer := 3840;
        YY19XX27        : integer := 3840;
        YY19XX28        : integer := 3840;
        YY20XX1         : integer := 1892;
        YY20XX2         : integer := 2985;
        YY20XX3         : integer := 3805;
        YY20XX4         : integer := 4078;
        YY20XX5         : integer := 3822;
        YY20XX6         : integer := 4095;
        YY20XX7         : integer := 4095;
        YY20XX8         : integer := 4095;
        YY20XX9         : integer := 4095;
        YY20XX10        : integer := 4095;
        YY20XX11        : integer := 4095;
        YY20XX12        : integer := 4095;
        YY20XX13        : integer := 4095;
        YY20XX14        : integer := 4095;
        YY20XX15        : integer := 4095;
        YY20XX16        : integer := 4095;
        YY20XX17        : integer := 4095;
        YY20XX18        : integer := 4095;
        YY20XX19        : integer := 4095;
        YY20XX20        : integer := 4095;
        YY20XX21        : integer := 4095;
        YY20XX22        : integer := 4095;
        YY20XX23        : integer := 4095;
        YY20XX24        : integer := 3565;
        YY20XX25        : integer := 1927;
        YY20XX26        : integer := 3840;
        YY20XX27        : integer := 3840;
        YY20XX28        : integer := 3840;
        YY21XX1         : integer := 2438;
        YY21XX2         : integer := 3258;
        YY21XX3         : integer := 4078;
        YY21XX4         : integer := 4095;
        YY21XX5         : integer := 4095;
        YY21XX6         : integer := 4095;
        YY21XX7         : integer := 4095;
        YY21XX8         : integer := 4095;
        YY21XX9         : integer := 4095;
        YY21XX10        : integer := 4095;
        YY21XX11        : integer := 4095;
        YY21XX12        : integer := 4095;
        YY21XX13        : integer := 4095;
        YY21XX14        : integer := 4095;
        YY21XX15        : integer := 4095;
        YY21XX16        : integer := 4095;
        YY21XX17        : integer := 4095;
        YY21XX18        : integer := 4095;
        YY21XX19        : integer := 4095;
        YY21XX20        : integer := 4095;
        YY21XX21        : integer := 4095;
        YY21XX22        : integer := 4095;
        YY21XX23        : integer := 4095;
        YY21XX24        : integer := 3276;
        YY21XX25        : integer := 1927;
        YY21XX26        : integer := 3840;
        YY21XX27        : integer := 3840;
        YY21XX28        : integer := 3840;
        YY22XX1         : integer := 2712;
        YY22XX2         : integer := 3531;
        YY22XX3         : integer := 4094;
        YY22XX4         : integer := 4095;
        YY22XX5         : integer := 4095;
        YY22XX6         : integer := 4095;
        YY22XX7         : integer := 4095;
        YY22XX8         : integer := 4095;
        YY22XX9         : integer := 4095;
        YY22XX10        : integer := 4095;
        YY22XX11        : integer := 4095;
        YY22XX12        : integer := 4095;
        YY22XX13        : integer := 4095;
        YY22XX14        : integer := 4095;
        YY22XX15        : integer := 4095;
        YY22XX16        : integer := 4095;
        YY22XX17        : integer := 4095;
        YY22XX18        : integer := 4095;
        YY22XX19        : integer := 4095;
        YY22XX20        : integer := 4095;
        YY22XX21        : integer := 4095;
        YY22XX22        : integer := 4095;
        YY22XX23        : integer := 3822;
        YY22XX24        : integer := 3276;
        YY22XX25        : integer := 2457;
        YY22XX26        : integer := 1911;
        YY22XX27        : integer := 1365;
        YY22XX28        : integer := 3840;
        YY23XX1         : integer := 2985;
        YY23XX2         : integer := 3548;
        YY23XX3         : integer := 4095;
        YY23XX4         : integer := 4095;
        YY23XX5         : integer := 4095;
        YY23XX6         : integer := 4095;
        YY23XX7         : integer := 4095;
        YY23XX8         : integer := 4095;
        YY23XX9         : integer := 4095;
        YY23XX10        : integer := 4095;
        YY23XX11        : integer := 4095;
        YY23XX12        : integer := 4095;
        YY23XX13        : integer := 4095;
        YY23XX14        : integer := 4095;
        YY23XX15        : integer := 4095;
        YY23XX16        : integer := 4095;
        YY23XX17        : integer := 4095;
        YY23XX18        : integer := 4095;
        YY23XX19        : integer := 4095;
        YY23XX20        : integer := 4095;
        YY23XX21        : integer := 4095;
        YY23XX22        : integer := 3822;
        YY23XX23        : integer := 3019;
        YY23XX24        : integer := 3003;
        YY23XX25        : integer := 3003;
        YY23XX26        : integer := 3276;
        YY23XX27        : integer := 3003;
        YY23XX28        : integer := 2183;
        YY24XX1         : integer := 2456;
        YY24XX2         : integer := 3019;
        YY24XX3         : integer := 3822;
        YY24XX4         : integer := 4095;
        YY24XX5         : integer := 4095;
        YY24XX6         : integer := 4095;
        YY24XX7         : integer := 4095;
        YY24XX8         : integer := 4095;
        YY24XX9         : integer := 4095;
        YY24XX10        : integer := 4095;
        YY24XX11        : integer := 4095;
        YY24XX12        : integer := 4095;
        YY24XX13        : integer := 4095;
        YY24XX14        : integer := 4095;
        YY24XX15        : integer := 4095;
        YY24XX16        : integer := 4095;
        YY24XX17        : integer := 4095;
        YY24XX18        : integer := 4095;
        YY24XX19        : integer := 4095;
        YY24XX20        : integer := 4095;
        YY24XX21        : integer := 4079;
        YY24XX22        : integer := 3822;
        YY24XX23        : integer := 3822;
        YY24XX24        : integer := 3566;
        YY24XX25        : integer := 3822;
        YY24XX26        : integer := 4095;
        YY24XX27        : integer := 3822;
        YY24XX28        : integer := 2729;
        YY25XX1         : integer := 1638;
        YY25XX2         : integer := 2184;
        YY25XX3         : integer := 3003;
        YY25XX4         : integer := 3566;
        YY25XX5         : integer := 3839;
        YY25XX6         : integer := 4095;
        YY25XX7         : integer := 4095;
        YY25XX8         : integer := 4095;
        YY25XX9         : integer := 4095;
        YY25XX10        : integer := 4095;
        YY25XX11        : integer := 4095;
        YY25XX12        : integer := 4095;
        YY25XX13        : integer := 4095;
        YY25XX14        : integer := 4095;
        YY25XX15        : integer := 4095;
        YY25XX16        : integer := 4095;
        YY25XX17        : integer := 4095;
        YY25XX18        : integer := 4095;
        YY25XX19        : integer := 4079;
        YY25XX20        : integer := 4078;
        YY25XX21        : integer := 4079;
        YY25XX22        : integer := 3822;
        YY25XX23        : integer := 4095;
        YY25XX24        : integer := 4095;
        YY25XX25        : integer := 4095;
        YY25XX26        : integer := 4095;
        YY25XX27        : integer := 3275;
        YY25XX28        : integer := 1910;
        YY26XX1         : integer := 819;
        YY26XX2         : integer := 1365;
        YY26XX3         : integer := 1928;
        YY26XX4         : integer := 3020;
        YY26XX5         : integer := 3294;
        YY26XX6         : integer := 3823;
        YY26XX7         : integer := 3823;
        YY26XX8         : integer := 4079;
        YY26XX9         : integer := 4095;
        YY26XX10        : integer := 4095;
        YY26XX11        : integer := 4095;
        YY26XX12        : integer := 4095;
        YY26XX13        : integer := 4095;
        YY26XX14        : integer := 4095;
        YY26XX15        : integer := 4095;
        YY26XX16        : integer := 4095;
        YY26XX17        : integer := 4095;
        YY26XX18        : integer := 3806;
        YY26XX19        : integer := 3549;
        YY26XX20        : integer := 3806;
        YY26XX21        : integer := 4079;
        YY26XX22        : integer := 4095;
        YY26XX23        : integer := 4095;
        YY26XX24        : integer := 4095;
        YY26XX25        : integer := 4095;
        YY26XX26        : integer := 3003;
        YY26XX27        : integer := 1910;
        YY26XX28        : integer := 819;
        YY27XX1         : integer := 3840;
        YY27XX2         : integer := 563;
        YY27XX3         : integer := 1109;
        YY27XX4         : integer := 1928;
        YY27XX5         : integer := 2474;
        YY27XX6         : integer := 3277;
        YY27XX7         : integer := 3549;
        YY27XX8         : integer := 3550;
        YY27XX9         : integer := 3806;
        YY27XX10        : integer := 3822;
        YY27XX11        : integer := 3823;
        YY27XX12        : integer := 4079;
        YY27XX13        : integer := 4079;
        YY27XX14        : integer := 4079;
        YY27XX15        : integer := 4079;
        YY27XX16        : integer := 3822;
        YY27XX17        : integer := 3549;
        YY27XX18        : integer := 3276;
        YY27XX19        : integer := 3276;
        YY27XX20        : integer := 3806;
        YY27XX21        : integer := 4095;
        YY27XX22        : integer := 4095;
        YY27XX23        : integer := 4095;
        YY27XX24        : integer := 4095;
        YY27XX25        : integer := 3003;
        YY27XX26        : integer := 1911;
        YY27XX27        : integer := 819;
        YY27XX28        : integer := 3840;
        YY28XX1         : integer := 3840;
        YY28XX2         : integer := 3840;
        YY28XX3         : integer := 546;
        YY28XX4         : integer := 1093;
        YY28XX5         : integer := 1639;
        YY28XX6         : integer := 2458;
        YY28XX7         : integer := 3004;
        YY28XX8         : integer := 3260;
        YY28XX9         : integer := 3276;
        YY28XX10        : integer := 3276;
        YY28XX11        : integer := 3533;
        YY28XX12        : integer := 3533;
        YY28XX13        : integer := 3533;
        YY28XX14        : integer := 3533;
        YY28XX15        : integer := 3533;
        YY28XX16        : integer := 3276;
        YY28XX17        : integer := 3003;
        YY28XX18        : integer := 3003;
        YY28XX19        : integer := 3276;
        YY28XX20        : integer := 4079;
        YY28XX21        : integer := 4095;
        YY28XX22        : integer := 4095;
        YY28XX23        : integer := 3822;
        YY28XX24        : integer := 3003;
        YY28XX25        : integer := 1638;
        YY28XX26        : integer := 546;
        YY28XX27        : integer := 3840;
        YY28XX28        : integer := 3840;
        YY29XX1         : integer := 3840;
        YY29XX2         : integer := 3840;
        YY29XX3         : integer := 3840;
        YY29XX4         : integer := 3840;
        YY29XX5         : integer := 1075;
        YY29XX6         : integer := 1365;
        YY29XX7         : integer := 2168;
        YY29XX8         : integer := 2440;
        YY29XX9         : integer := 2457;
        YY29XX10        : integer := 2457;
        YY29XX11        : integer := 2457;
        YY29XX12        : integer := 2458;
        YY29XX13        : integer := 2714;
        YY29XX14        : integer := 2457;
        YY29XX15        : integer := 2184;
        YY29XX16        : integer := 2457;
        YY29XX17        : integer := 2714;
        YY29XX18        : integer := 3003;
        YY29XX19        : integer := 3550;
        YY29XX20        : integer := 4095;
        YY29XX21        : integer := 4095;
        YY29XX22        : integer := 3549;
        YY29XX23        : integer := 2184;
        YY29XX24        : integer := 1364;
        YY29XX25        : integer := 273;
        YY29XX26        : integer := 3840;
        YY29XX27        : integer := 3840;
        YY29XX28        : integer := 3840;
        YY30XX1         : integer := 3840;
        YY30XX2         : integer := 3840;
        YY30XX3         : integer := 3840;
        YY30XX4         : integer := 3840;
        YY30XX5         : integer := 3840;
        YY30XX6         : integer := 802;
        YY30XX7         : integer := 1092;
        YY30XX8         : integer := 1365;
        YY30XX9         : integer := 1638;
        YY30XX10        : integer := 1911;
        YY30XX11        : integer := 1911;
        YY30XX12        : integer := 1638;
        YY30XX13        : integer := 1638;
        YY30XX14        : integer := 1895;
        YY30XX15        : integer := 1895;
        YY30XX16        : integer := 1911;
        YY30XX17        : integer := 2441;
        YY30XX18        : integer := 2987;
        YY30XX19        : integer := 3549;
        YY30XX20        : integer := 3822;
        YY30XX21        : integer := 3003;
        YY30XX22        : integer := 1911;
        YY30XX23        : integer := 1348;
        YY30XX24        : integer := 818;
        YY30XX25        : integer := 3840;
        YY30XX26        : integer := 3840;
        YY30XX27        : integer := 3840;
        YY30XX28        : integer := 3840;
        YY31XX1         : integer := 3840;
        YY31XX2         : integer := 3840;
        YY31XX3         : integer := 3840;
        YY31XX4         : integer := 3840;
        YY31XX5         : integer := 3840;
        YY31XX6         : integer := 3840;
        YY31XX7         : integer := 3840;
        YY31XX8         : integer := 819;
        YY31XX9         : integer := 1348;
        YY31XX10        : integer := 1638;
        YY31XX11        : integer := 1365;
        YY31XX12        : integer := 1348;
        YY31XX13        : integer := 1365;
        YY31XX14        : integer := 1638;
        YY31XX15        : integer := 1895;
        YY31XX16        : integer := 2184;
        YY31XX17        : integer := 2457;
        YY31XX18        : integer := 2987;
        YY31XX19        : integer := 3276;
        YY31XX20        : integer := 3003;
        YY31XX21        : integer := 1911;
        YY31XX22        : integer := 803;
        YY31XX23        : integer := 546;
        YY31XX24        : integer := 3840;
        YY31XX25        : integer := 3840;
        YY31XX26        : integer := 3840;
        YY31XX27        : integer := 3840;
        YY31XX28        : integer := 3840;
        YY32XX1         : integer := 3840;
        YY32XX2         : integer := 3840;
        YY32XX3         : integer := 3840;
        YY32XX4         : integer := 3840;
        YY32XX5         : integer := 3840;
        YY32XX6         : integer := 3840;
        YY32XX7         : integer := 3840;
        YY32XX8         : integer := 3840;
        YY32XX9         : integer := 3840;
        YY32XX10        : integer := 3840;
        YY32XX11        : integer := 3840;
        YY32XX12        : integer := 3840;
        YY32XX13        : integer := 3840;
        YY32XX14        : integer := 1365;
        YY32XX15        : integer := 2167;
        YY32XX16        : integer := 2713;
        YY32XX17        : integer := 2986;
        YY32XX18        : integer := 2714;
        YY32XX19        : integer := 2168;
        YY32XX20        : integer := 1622;
        YY32XX21        : integer := 1076;
        YY32XX22        : integer := 546;
        YY32XX23        : integer := 3840;
        YY32XX24        : integer := 3840;
        YY32XX25        : integer := 3840;
        YY32XX26        : integer := 3840;
        YY32XX27        : integer := 3840;
        YY32XX28        : integer := 3840;
        YY33XX1         : integer := 3840;
        YY33XX2         : integer := 3840;
        YY33XX3         : integer := 3840;
        YY33XX4         : integer := 3840;
        YY33XX5         : integer := 3840;
        YY33XX6         : integer := 3840;
        YY33XX7         : integer := 3840;
        YY33XX8         : integer := 3840;
        YY33XX9         : integer := 3840;
        YY33XX10        : integer := 3840;
        YY33XX11        : integer := 3840;
        YY33XX12        : integer := 3840;
        YY33XX13        : integer := 3840;
        YY33XX14        : integer := 1091;
        YY33XX15        : integer := 1910;
        YY33XX16        : integer := 2184;
        YY33XX17        : integer := 2184;
        YY33XX18        : integer := 1638;
        YY33XX19        : integer := 819;
        YY33XX20        : integer := 546;
        YY33XX21        : integer := 546;
        YY33XX22        : integer := 3840;
        YY33XX23        : integer := 3840;
        YY33XX24        : integer := 3840;
        YY33XX25        : integer := 3840;
        YY33XX26        : integer := 3840;
        YY33XX27        : integer := 3840;
        YY33XX28        : integer := 3840;
        YY34XX1         : integer := 3840;
        YY34XX2         : integer := 3840;
        YY34XX3         : integer := 3840;
        YY34XX4         : integer := 3840;
        YY34XX5         : integer := 3840;
        YY34XX6         : integer := 3840;
        YY34XX7         : integer := 3840;
        YY34XX8         : integer := 3840;
        YY34XX9         : integer := 3840;
        YY34XX10        : integer := 3840;
        YY34XX11        : integer := 3840;
        YY34XX12        : integer := 3840;
        YY34XX13        : integer := 3840;
        YY34XX14        : integer := 818;
        YY34XX15        : integer := 1348;
        YY34XX16        : integer := 1364;
        YY34XX17        : integer := 1092;
        YY34XX18        : integer := 819;
        YY34XX19        : integer := 546;
        YY34XX20        : integer := 3840;
        YY34XX21        : integer := 3840;
        YY34XX22        : integer := 3840;
        YY34XX23        : integer := 3840;
        YY34XX24        : integer := 3840;
        YY34XX25        : integer := 3840;
        YY34XX26        : integer := 3840;
        YY34XX27        : integer := 3840;
        YY34XX28        : integer := 3840;
        YY35XX1         : integer := 3840;
        YY35XX2         : integer := 3840;
        YY35XX3         : integer := 3840;
        YY35XX4         : integer := 3840;
        YY35XX5         : integer := 3840;
        YY35XX6         : integer := 3840;
        YY35XX7         : integer := 3840;
        YY35XX8         : integer := 3840;
        YY35XX9         : integer := 3840;
        YY35XX10        : integer := 3840;
        YY35XX11        : integer := 3840;
        YY35XX12        : integer := 3840;
        YY35XX13        : integer := 3840;
        YY35XX14        : integer := 3840;
        YY35XX15        : integer := 818;
        YY35XX16        : integer := 802;
        YY35XX17        : integer := 546;
        YY35XX18        : integer := 545;
        YY35XX19        : integer := 3840;
        YY35XX20        : integer := 3840;
        YY35XX21        : integer := 3840;
        YY35XX22        : integer := 3840;
        YY35XX23        : integer := 3840;
        YY35XX24        : integer := 3840;
        YY35XX25        : integer := 3840;
        YY35XX26        : integer := 3840;
        YY35XX27        : integer := 3840;
        YY35XX28        : integer := 3840
    );
    port(
        RGB             : out    vl_logic_vector(11 downto 0);
        YX              : in     vl_logic_vector(19 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of Y0X0 : constant is 1;
    attribute mti_svvh_generic_type of Y0X1 : constant is 1;
    attribute mti_svvh_generic_type of Y0X2 : constant is 1;
    attribute mti_svvh_generic_type of Y0X3 : constant is 1;
    attribute mti_svvh_generic_type of Y0X4 : constant is 1;
    attribute mti_svvh_generic_type of Y0X5 : constant is 1;
    attribute mti_svvh_generic_type of Y0X6 : constant is 1;
    attribute mti_svvh_generic_type of Y0X7 : constant is 1;
    attribute mti_svvh_generic_type of Y0X8 : constant is 1;
    attribute mti_svvh_generic_type of Y0X9 : constant is 1;
    attribute mti_svvh_generic_type of Y0X10 : constant is 1;
    attribute mti_svvh_generic_type of Y0X11 : constant is 1;
    attribute mti_svvh_generic_type of Y0X12 : constant is 1;
    attribute mti_svvh_generic_type of Y0X13 : constant is 1;
    attribute mti_svvh_generic_type of Y0X14 : constant is 1;
    attribute mti_svvh_generic_type of Y0X15 : constant is 1;
    attribute mti_svvh_generic_type of Y0X16 : constant is 1;
    attribute mti_svvh_generic_type of Y0X17 : constant is 1;
    attribute mti_svvh_generic_type of Y0X18 : constant is 1;
    attribute mti_svvh_generic_type of Y0X19 : constant is 1;
    attribute mti_svvh_generic_type of Y0X20 : constant is 1;
    attribute mti_svvh_generic_type of Y0X21 : constant is 1;
    attribute mti_svvh_generic_type of Y0X22 : constant is 1;
    attribute mti_svvh_generic_type of Y0X23 : constant is 1;
    attribute mti_svvh_generic_type of Y0X24 : constant is 1;
    attribute mti_svvh_generic_type of Y0X25 : constant is 1;
    attribute mti_svvh_generic_type of Y0X26 : constant is 1;
    attribute mti_svvh_generic_type of Y0X27 : constant is 1;
    attribute mti_svvh_generic_type of Y0X28 : constant is 1;
    attribute mti_svvh_generic_type of Y1X1 : constant is 1;
    attribute mti_svvh_generic_type of Y1X2 : constant is 1;
    attribute mti_svvh_generic_type of Y1X3 : constant is 1;
    attribute mti_svvh_generic_type of Y1X4 : constant is 1;
    attribute mti_svvh_generic_type of Y1X5 : constant is 1;
    attribute mti_svvh_generic_type of Y1X6 : constant is 1;
    attribute mti_svvh_generic_type of Y1X7 : constant is 1;
    attribute mti_svvh_generic_type of Y1X8 : constant is 1;
    attribute mti_svvh_generic_type of Y1X9 : constant is 1;
    attribute mti_svvh_generic_type of Y1X10 : constant is 1;
    attribute mti_svvh_generic_type of Y1X11 : constant is 1;
    attribute mti_svvh_generic_type of Y1X12 : constant is 1;
    attribute mti_svvh_generic_type of Y1X13 : constant is 1;
    attribute mti_svvh_generic_type of Y1X14 : constant is 1;
    attribute mti_svvh_generic_type of Y1X15 : constant is 1;
    attribute mti_svvh_generic_type of Y1X16 : constant is 1;
    attribute mti_svvh_generic_type of Y1X17 : constant is 1;
    attribute mti_svvh_generic_type of Y1X18 : constant is 1;
    attribute mti_svvh_generic_type of Y1X19 : constant is 1;
    attribute mti_svvh_generic_type of Y1X20 : constant is 1;
    attribute mti_svvh_generic_type of Y1X21 : constant is 1;
    attribute mti_svvh_generic_type of Y1X22 : constant is 1;
    attribute mti_svvh_generic_type of Y1X23 : constant is 1;
    attribute mti_svvh_generic_type of Y1X24 : constant is 1;
    attribute mti_svvh_generic_type of Y1X25 : constant is 1;
    attribute mti_svvh_generic_type of Y1X26 : constant is 1;
    attribute mti_svvh_generic_type of Y1X27 : constant is 1;
    attribute mti_svvh_generic_type of Y1X28 : constant is 1;
    attribute mti_svvh_generic_type of Y2X1 : constant is 1;
    attribute mti_svvh_generic_type of Y2X2 : constant is 1;
    attribute mti_svvh_generic_type of Y2X3 : constant is 1;
    attribute mti_svvh_generic_type of Y2X4 : constant is 1;
    attribute mti_svvh_generic_type of Y2X5 : constant is 1;
    attribute mti_svvh_generic_type of Y2X6 : constant is 1;
    attribute mti_svvh_generic_type of Y2X7 : constant is 1;
    attribute mti_svvh_generic_type of Y2X8 : constant is 1;
    attribute mti_svvh_generic_type of Y2X9 : constant is 1;
    attribute mti_svvh_generic_type of Y2X10 : constant is 1;
    attribute mti_svvh_generic_type of Y2X11 : constant is 1;
    attribute mti_svvh_generic_type of Y2X12 : constant is 1;
    attribute mti_svvh_generic_type of Y2X13 : constant is 1;
    attribute mti_svvh_generic_type of Y2X14 : constant is 1;
    attribute mti_svvh_generic_type of Y2X15 : constant is 1;
    attribute mti_svvh_generic_type of Y2X16 : constant is 1;
    attribute mti_svvh_generic_type of Y2X17 : constant is 1;
    attribute mti_svvh_generic_type of Y2X18 : constant is 1;
    attribute mti_svvh_generic_type of Y2X19 : constant is 1;
    attribute mti_svvh_generic_type of Y2X20 : constant is 1;
    attribute mti_svvh_generic_type of Y2X21 : constant is 1;
    attribute mti_svvh_generic_type of Y2X22 : constant is 1;
    attribute mti_svvh_generic_type of Y2X23 : constant is 1;
    attribute mti_svvh_generic_type of Y2X24 : constant is 1;
    attribute mti_svvh_generic_type of Y2X25 : constant is 1;
    attribute mti_svvh_generic_type of Y2X26 : constant is 1;
    attribute mti_svvh_generic_type of Y2X27 : constant is 1;
    attribute mti_svvh_generic_type of Y2X28 : constant is 1;
    attribute mti_svvh_generic_type of Y3X1 : constant is 1;
    attribute mti_svvh_generic_type of Y3X2 : constant is 1;
    attribute mti_svvh_generic_type of Y3X3 : constant is 1;
    attribute mti_svvh_generic_type of Y3X4 : constant is 1;
    attribute mti_svvh_generic_type of Y3X5 : constant is 1;
    attribute mti_svvh_generic_type of Y3X6 : constant is 1;
    attribute mti_svvh_generic_type of Y3X7 : constant is 1;
    attribute mti_svvh_generic_type of Y3X8 : constant is 1;
    attribute mti_svvh_generic_type of Y3X9 : constant is 1;
    attribute mti_svvh_generic_type of Y3X10 : constant is 1;
    attribute mti_svvh_generic_type of Y3X11 : constant is 1;
    attribute mti_svvh_generic_type of Y3X12 : constant is 1;
    attribute mti_svvh_generic_type of Y3X13 : constant is 1;
    attribute mti_svvh_generic_type of Y3X14 : constant is 1;
    attribute mti_svvh_generic_type of Y3X15 : constant is 1;
    attribute mti_svvh_generic_type of Y3X16 : constant is 1;
    attribute mti_svvh_generic_type of Y3X17 : constant is 1;
    attribute mti_svvh_generic_type of Y3X18 : constant is 1;
    attribute mti_svvh_generic_type of Y3X19 : constant is 1;
    attribute mti_svvh_generic_type of Y3X20 : constant is 1;
    attribute mti_svvh_generic_type of Y3X21 : constant is 1;
    attribute mti_svvh_generic_type of Y3X22 : constant is 1;
    attribute mti_svvh_generic_type of Y3X23 : constant is 1;
    attribute mti_svvh_generic_type of Y3X24 : constant is 1;
    attribute mti_svvh_generic_type of Y3X25 : constant is 1;
    attribute mti_svvh_generic_type of Y3X26 : constant is 1;
    attribute mti_svvh_generic_type of Y3X27 : constant is 1;
    attribute mti_svvh_generic_type of Y3X28 : constant is 1;
    attribute mti_svvh_generic_type of Y4X1 : constant is 1;
    attribute mti_svvh_generic_type of Y4X2 : constant is 1;
    attribute mti_svvh_generic_type of Y4X3 : constant is 1;
    attribute mti_svvh_generic_type of Y4X4 : constant is 1;
    attribute mti_svvh_generic_type of Y4X5 : constant is 1;
    attribute mti_svvh_generic_type of Y4X6 : constant is 1;
    attribute mti_svvh_generic_type of Y4X7 : constant is 1;
    attribute mti_svvh_generic_type of Y4X8 : constant is 1;
    attribute mti_svvh_generic_type of Y4X9 : constant is 1;
    attribute mti_svvh_generic_type of Y4X10 : constant is 1;
    attribute mti_svvh_generic_type of Y4X11 : constant is 1;
    attribute mti_svvh_generic_type of Y4X12 : constant is 1;
    attribute mti_svvh_generic_type of Y4X13 : constant is 1;
    attribute mti_svvh_generic_type of Y4X14 : constant is 1;
    attribute mti_svvh_generic_type of Y4X15 : constant is 1;
    attribute mti_svvh_generic_type of Y4X16 : constant is 1;
    attribute mti_svvh_generic_type of Y4X17 : constant is 1;
    attribute mti_svvh_generic_type of Y4X18 : constant is 1;
    attribute mti_svvh_generic_type of Y4X19 : constant is 1;
    attribute mti_svvh_generic_type of Y4X20 : constant is 1;
    attribute mti_svvh_generic_type of Y4X21 : constant is 1;
    attribute mti_svvh_generic_type of Y4X22 : constant is 1;
    attribute mti_svvh_generic_type of Y4X23 : constant is 1;
    attribute mti_svvh_generic_type of Y4X24 : constant is 1;
    attribute mti_svvh_generic_type of Y4X25 : constant is 1;
    attribute mti_svvh_generic_type of Y4X26 : constant is 1;
    attribute mti_svvh_generic_type of Y4X27 : constant is 1;
    attribute mti_svvh_generic_type of Y4X28 : constant is 1;
    attribute mti_svvh_generic_type of Y5X1 : constant is 1;
    attribute mti_svvh_generic_type of Y5X2 : constant is 1;
    attribute mti_svvh_generic_type of Y5X3 : constant is 1;
    attribute mti_svvh_generic_type of Y5X4 : constant is 1;
    attribute mti_svvh_generic_type of Y5X5 : constant is 1;
    attribute mti_svvh_generic_type of Y5X6 : constant is 1;
    attribute mti_svvh_generic_type of Y5X7 : constant is 1;
    attribute mti_svvh_generic_type of Y5X8 : constant is 1;
    attribute mti_svvh_generic_type of Y5X9 : constant is 1;
    attribute mti_svvh_generic_type of Y5X10 : constant is 1;
    attribute mti_svvh_generic_type of Y5X11 : constant is 1;
    attribute mti_svvh_generic_type of Y5X12 : constant is 1;
    attribute mti_svvh_generic_type of Y5X13 : constant is 1;
    attribute mti_svvh_generic_type of Y5X14 : constant is 1;
    attribute mti_svvh_generic_type of Y5X15 : constant is 1;
    attribute mti_svvh_generic_type of Y5X16 : constant is 1;
    attribute mti_svvh_generic_type of Y5X17 : constant is 1;
    attribute mti_svvh_generic_type of Y5X18 : constant is 1;
    attribute mti_svvh_generic_type of Y5X19 : constant is 1;
    attribute mti_svvh_generic_type of Y5X20 : constant is 1;
    attribute mti_svvh_generic_type of Y5X21 : constant is 1;
    attribute mti_svvh_generic_type of Y5X22 : constant is 1;
    attribute mti_svvh_generic_type of Y5X23 : constant is 1;
    attribute mti_svvh_generic_type of Y5X24 : constant is 1;
    attribute mti_svvh_generic_type of Y5X25 : constant is 1;
    attribute mti_svvh_generic_type of Y5X26 : constant is 1;
    attribute mti_svvh_generic_type of Y5X27 : constant is 1;
    attribute mti_svvh_generic_type of Y5X28 : constant is 1;
    attribute mti_svvh_generic_type of Y6X1 : constant is 1;
    attribute mti_svvh_generic_type of Y6X2 : constant is 1;
    attribute mti_svvh_generic_type of Y6X3 : constant is 1;
    attribute mti_svvh_generic_type of Y6X4 : constant is 1;
    attribute mti_svvh_generic_type of Y6X5 : constant is 1;
    attribute mti_svvh_generic_type of Y6X6 : constant is 1;
    attribute mti_svvh_generic_type of Y6X7 : constant is 1;
    attribute mti_svvh_generic_type of Y6X8 : constant is 1;
    attribute mti_svvh_generic_type of Y6X9 : constant is 1;
    attribute mti_svvh_generic_type of Y6X10 : constant is 1;
    attribute mti_svvh_generic_type of Y6X11 : constant is 1;
    attribute mti_svvh_generic_type of Y6X12 : constant is 1;
    attribute mti_svvh_generic_type of Y6X13 : constant is 1;
    attribute mti_svvh_generic_type of Y6X14 : constant is 1;
    attribute mti_svvh_generic_type of Y6X15 : constant is 1;
    attribute mti_svvh_generic_type of Y6X16 : constant is 1;
    attribute mti_svvh_generic_type of Y6X17 : constant is 1;
    attribute mti_svvh_generic_type of Y6X18 : constant is 1;
    attribute mti_svvh_generic_type of Y6X19 : constant is 1;
    attribute mti_svvh_generic_type of Y6X20 : constant is 1;
    attribute mti_svvh_generic_type of Y6X21 : constant is 1;
    attribute mti_svvh_generic_type of Y6X22 : constant is 1;
    attribute mti_svvh_generic_type of Y6X23 : constant is 1;
    attribute mti_svvh_generic_type of Y6X24 : constant is 1;
    attribute mti_svvh_generic_type of Y6X25 : constant is 1;
    attribute mti_svvh_generic_type of Y6X26 : constant is 1;
    attribute mti_svvh_generic_type of Y6X27 : constant is 1;
    attribute mti_svvh_generic_type of Y6X28 : constant is 1;
    attribute mti_svvh_generic_type of Y7X1 : constant is 1;
    attribute mti_svvh_generic_type of Y7X2 : constant is 1;
    attribute mti_svvh_generic_type of Y7X3 : constant is 1;
    attribute mti_svvh_generic_type of Y7X4 : constant is 1;
    attribute mti_svvh_generic_type of Y7X5 : constant is 1;
    attribute mti_svvh_generic_type of Y7X6 : constant is 1;
    attribute mti_svvh_generic_type of Y7X7 : constant is 1;
    attribute mti_svvh_generic_type of Y7X8 : constant is 1;
    attribute mti_svvh_generic_type of Y7X9 : constant is 1;
    attribute mti_svvh_generic_type of Y7X10 : constant is 1;
    attribute mti_svvh_generic_type of Y7X11 : constant is 1;
    attribute mti_svvh_generic_type of Y7X12 : constant is 1;
    attribute mti_svvh_generic_type of Y7X13 : constant is 1;
    attribute mti_svvh_generic_type of Y7X14 : constant is 1;
    attribute mti_svvh_generic_type of Y7X15 : constant is 1;
    attribute mti_svvh_generic_type of Y7X16 : constant is 1;
    attribute mti_svvh_generic_type of Y7X17 : constant is 1;
    attribute mti_svvh_generic_type of Y7X18 : constant is 1;
    attribute mti_svvh_generic_type of Y7X19 : constant is 1;
    attribute mti_svvh_generic_type of Y7X20 : constant is 1;
    attribute mti_svvh_generic_type of Y7X21 : constant is 1;
    attribute mti_svvh_generic_type of Y7X22 : constant is 1;
    attribute mti_svvh_generic_type of Y7X23 : constant is 1;
    attribute mti_svvh_generic_type of Y7X24 : constant is 1;
    attribute mti_svvh_generic_type of Y7X25 : constant is 1;
    attribute mti_svvh_generic_type of Y7X26 : constant is 1;
    attribute mti_svvh_generic_type of Y7X27 : constant is 1;
    attribute mti_svvh_generic_type of Y7X28 : constant is 1;
    attribute mti_svvh_generic_type of Y8X1 : constant is 1;
    attribute mti_svvh_generic_type of Y8X2 : constant is 1;
    attribute mti_svvh_generic_type of Y8X3 : constant is 1;
    attribute mti_svvh_generic_type of Y8X4 : constant is 1;
    attribute mti_svvh_generic_type of Y8X5 : constant is 1;
    attribute mti_svvh_generic_type of Y8X6 : constant is 1;
    attribute mti_svvh_generic_type of Y8X7 : constant is 1;
    attribute mti_svvh_generic_type of Y8X8 : constant is 1;
    attribute mti_svvh_generic_type of Y8X9 : constant is 1;
    attribute mti_svvh_generic_type of Y8X10 : constant is 1;
    attribute mti_svvh_generic_type of Y8X11 : constant is 1;
    attribute mti_svvh_generic_type of Y8X12 : constant is 1;
    attribute mti_svvh_generic_type of Y8X13 : constant is 1;
    attribute mti_svvh_generic_type of Y8X14 : constant is 1;
    attribute mti_svvh_generic_type of Y8X15 : constant is 1;
    attribute mti_svvh_generic_type of Y8X16 : constant is 1;
    attribute mti_svvh_generic_type of Y8X17 : constant is 1;
    attribute mti_svvh_generic_type of Y8X18 : constant is 1;
    attribute mti_svvh_generic_type of Y8X19 : constant is 1;
    attribute mti_svvh_generic_type of Y8X20 : constant is 1;
    attribute mti_svvh_generic_type of Y8X21 : constant is 1;
    attribute mti_svvh_generic_type of Y8X22 : constant is 1;
    attribute mti_svvh_generic_type of Y8X23 : constant is 1;
    attribute mti_svvh_generic_type of Y8X24 : constant is 1;
    attribute mti_svvh_generic_type of Y8X25 : constant is 1;
    attribute mti_svvh_generic_type of Y8X26 : constant is 1;
    attribute mti_svvh_generic_type of Y8X27 : constant is 1;
    attribute mti_svvh_generic_type of Y8X28 : constant is 1;
    attribute mti_svvh_generic_type of Y9X1 : constant is 1;
    attribute mti_svvh_generic_type of Y9X2 : constant is 1;
    attribute mti_svvh_generic_type of Y9X3 : constant is 1;
    attribute mti_svvh_generic_type of Y9X4 : constant is 1;
    attribute mti_svvh_generic_type of Y9X5 : constant is 1;
    attribute mti_svvh_generic_type of Y9X6 : constant is 1;
    attribute mti_svvh_generic_type of Y9X7 : constant is 1;
    attribute mti_svvh_generic_type of Y9X8 : constant is 1;
    attribute mti_svvh_generic_type of Y9X9 : constant is 1;
    attribute mti_svvh_generic_type of Y9X10 : constant is 1;
    attribute mti_svvh_generic_type of Y9X11 : constant is 1;
    attribute mti_svvh_generic_type of Y9X12 : constant is 1;
    attribute mti_svvh_generic_type of Y9X13 : constant is 1;
    attribute mti_svvh_generic_type of Y9X14 : constant is 1;
    attribute mti_svvh_generic_type of Y9X15 : constant is 1;
    attribute mti_svvh_generic_type of Y9X16 : constant is 1;
    attribute mti_svvh_generic_type of Y9X17 : constant is 1;
    attribute mti_svvh_generic_type of Y9X18 : constant is 1;
    attribute mti_svvh_generic_type of Y9X19 : constant is 1;
    attribute mti_svvh_generic_type of Y9X20 : constant is 1;
    attribute mti_svvh_generic_type of Y9X21 : constant is 1;
    attribute mti_svvh_generic_type of Y9X22 : constant is 1;
    attribute mti_svvh_generic_type of Y9X23 : constant is 1;
    attribute mti_svvh_generic_type of Y9X24 : constant is 1;
    attribute mti_svvh_generic_type of Y9X25 : constant is 1;
    attribute mti_svvh_generic_type of Y9X26 : constant is 1;
    attribute mti_svvh_generic_type of Y9X27 : constant is 1;
    attribute mti_svvh_generic_type of Y9X28 : constant is 1;
    attribute mti_svvh_generic_type of Y10X1 : constant is 1;
    attribute mti_svvh_generic_type of Y10X2 : constant is 1;
    attribute mti_svvh_generic_type of Y10X3 : constant is 1;
    attribute mti_svvh_generic_type of Y10X4 : constant is 1;
    attribute mti_svvh_generic_type of Y10X5 : constant is 1;
    attribute mti_svvh_generic_type of Y10X6 : constant is 1;
    attribute mti_svvh_generic_type of Y10X7 : constant is 1;
    attribute mti_svvh_generic_type of Y10X8 : constant is 1;
    attribute mti_svvh_generic_type of Y10X9 : constant is 1;
    attribute mti_svvh_generic_type of Y10X10 : constant is 1;
    attribute mti_svvh_generic_type of Y10X11 : constant is 1;
    attribute mti_svvh_generic_type of Y10X12 : constant is 1;
    attribute mti_svvh_generic_type of Y10X13 : constant is 1;
    attribute mti_svvh_generic_type of Y10X14 : constant is 1;
    attribute mti_svvh_generic_type of Y10X15 : constant is 1;
    attribute mti_svvh_generic_type of Y10X16 : constant is 1;
    attribute mti_svvh_generic_type of Y10X17 : constant is 1;
    attribute mti_svvh_generic_type of Y10X18 : constant is 1;
    attribute mti_svvh_generic_type of Y10X19 : constant is 1;
    attribute mti_svvh_generic_type of Y10X20 : constant is 1;
    attribute mti_svvh_generic_type of Y10X21 : constant is 1;
    attribute mti_svvh_generic_type of Y10X22 : constant is 1;
    attribute mti_svvh_generic_type of Y10X23 : constant is 1;
    attribute mti_svvh_generic_type of Y10X24 : constant is 1;
    attribute mti_svvh_generic_type of Y10X25 : constant is 1;
    attribute mti_svvh_generic_type of Y10X26 : constant is 1;
    attribute mti_svvh_generic_type of Y10X27 : constant is 1;
    attribute mti_svvh_generic_type of Y10X28 : constant is 1;
    attribute mti_svvh_generic_type of Y11X1 : constant is 1;
    attribute mti_svvh_generic_type of Y11X2 : constant is 1;
    attribute mti_svvh_generic_type of Y11X3 : constant is 1;
    attribute mti_svvh_generic_type of Y11X4 : constant is 1;
    attribute mti_svvh_generic_type of Y11X5 : constant is 1;
    attribute mti_svvh_generic_type of Y11X6 : constant is 1;
    attribute mti_svvh_generic_type of Y11X7 : constant is 1;
    attribute mti_svvh_generic_type of Y11X8 : constant is 1;
    attribute mti_svvh_generic_type of Y11X9 : constant is 1;
    attribute mti_svvh_generic_type of Y11X10 : constant is 1;
    attribute mti_svvh_generic_type of Y11X11 : constant is 1;
    attribute mti_svvh_generic_type of Y11X12 : constant is 1;
    attribute mti_svvh_generic_type of Y11X13 : constant is 1;
    attribute mti_svvh_generic_type of Y11X14 : constant is 1;
    attribute mti_svvh_generic_type of Y11X15 : constant is 1;
    attribute mti_svvh_generic_type of Y11X16 : constant is 1;
    attribute mti_svvh_generic_type of Y11X17 : constant is 1;
    attribute mti_svvh_generic_type of Y11X18 : constant is 1;
    attribute mti_svvh_generic_type of Y11X19 : constant is 1;
    attribute mti_svvh_generic_type of Y11X20 : constant is 1;
    attribute mti_svvh_generic_type of Y11X21 : constant is 1;
    attribute mti_svvh_generic_type of Y11X22 : constant is 1;
    attribute mti_svvh_generic_type of Y11X23 : constant is 1;
    attribute mti_svvh_generic_type of Y11X24 : constant is 1;
    attribute mti_svvh_generic_type of Y11X25 : constant is 1;
    attribute mti_svvh_generic_type of Y11X26 : constant is 1;
    attribute mti_svvh_generic_type of Y11X27 : constant is 1;
    attribute mti_svvh_generic_type of Y11X28 : constant is 1;
    attribute mti_svvh_generic_type of Y12X1 : constant is 1;
    attribute mti_svvh_generic_type of Y12X2 : constant is 1;
    attribute mti_svvh_generic_type of Y12X3 : constant is 1;
    attribute mti_svvh_generic_type of Y12X4 : constant is 1;
    attribute mti_svvh_generic_type of Y12X5 : constant is 1;
    attribute mti_svvh_generic_type of Y12X6 : constant is 1;
    attribute mti_svvh_generic_type of Y12X7 : constant is 1;
    attribute mti_svvh_generic_type of Y12X8 : constant is 1;
    attribute mti_svvh_generic_type of Y12X9 : constant is 1;
    attribute mti_svvh_generic_type of Y12X10 : constant is 1;
    attribute mti_svvh_generic_type of Y12X11 : constant is 1;
    attribute mti_svvh_generic_type of Y12X12 : constant is 1;
    attribute mti_svvh_generic_type of Y12X13 : constant is 1;
    attribute mti_svvh_generic_type of Y12X14 : constant is 1;
    attribute mti_svvh_generic_type of Y12X15 : constant is 1;
    attribute mti_svvh_generic_type of Y12X16 : constant is 1;
    attribute mti_svvh_generic_type of Y12X17 : constant is 1;
    attribute mti_svvh_generic_type of Y12X18 : constant is 1;
    attribute mti_svvh_generic_type of Y12X19 : constant is 1;
    attribute mti_svvh_generic_type of Y12X20 : constant is 1;
    attribute mti_svvh_generic_type of Y12X21 : constant is 1;
    attribute mti_svvh_generic_type of Y12X22 : constant is 1;
    attribute mti_svvh_generic_type of Y12X23 : constant is 1;
    attribute mti_svvh_generic_type of Y12X24 : constant is 1;
    attribute mti_svvh_generic_type of Y12X25 : constant is 1;
    attribute mti_svvh_generic_type of Y12X26 : constant is 1;
    attribute mti_svvh_generic_type of Y12X27 : constant is 1;
    attribute mti_svvh_generic_type of Y12X28 : constant is 1;
    attribute mti_svvh_generic_type of Y13X1 : constant is 1;
    attribute mti_svvh_generic_type of Y13X2 : constant is 1;
    attribute mti_svvh_generic_type of Y13X3 : constant is 1;
    attribute mti_svvh_generic_type of Y13X4 : constant is 1;
    attribute mti_svvh_generic_type of Y13X5 : constant is 1;
    attribute mti_svvh_generic_type of Y13X6 : constant is 1;
    attribute mti_svvh_generic_type of Y13X7 : constant is 1;
    attribute mti_svvh_generic_type of Y13X8 : constant is 1;
    attribute mti_svvh_generic_type of Y13X9 : constant is 1;
    attribute mti_svvh_generic_type of Y13X10 : constant is 1;
    attribute mti_svvh_generic_type of Y13X11 : constant is 1;
    attribute mti_svvh_generic_type of Y13X12 : constant is 1;
    attribute mti_svvh_generic_type of Y13X13 : constant is 1;
    attribute mti_svvh_generic_type of Y13X14 : constant is 1;
    attribute mti_svvh_generic_type of Y13X15 : constant is 1;
    attribute mti_svvh_generic_type of Y13X16 : constant is 1;
    attribute mti_svvh_generic_type of Y13X17 : constant is 1;
    attribute mti_svvh_generic_type of Y13X18 : constant is 1;
    attribute mti_svvh_generic_type of Y13X19 : constant is 1;
    attribute mti_svvh_generic_type of Y13X20 : constant is 1;
    attribute mti_svvh_generic_type of Y13X21 : constant is 1;
    attribute mti_svvh_generic_type of Y13X22 : constant is 1;
    attribute mti_svvh_generic_type of Y13X23 : constant is 1;
    attribute mti_svvh_generic_type of Y13X24 : constant is 1;
    attribute mti_svvh_generic_type of Y13X25 : constant is 1;
    attribute mti_svvh_generic_type of Y13X26 : constant is 1;
    attribute mti_svvh_generic_type of Y13X27 : constant is 1;
    attribute mti_svvh_generic_type of Y13X28 : constant is 1;
    attribute mti_svvh_generic_type of Y14X1 : constant is 1;
    attribute mti_svvh_generic_type of Y14X2 : constant is 1;
    attribute mti_svvh_generic_type of Y14X3 : constant is 1;
    attribute mti_svvh_generic_type of Y14X4 : constant is 1;
    attribute mti_svvh_generic_type of Y14X5 : constant is 1;
    attribute mti_svvh_generic_type of Y14X6 : constant is 1;
    attribute mti_svvh_generic_type of Y14X7 : constant is 1;
    attribute mti_svvh_generic_type of Y14X8 : constant is 1;
    attribute mti_svvh_generic_type of Y14X9 : constant is 1;
    attribute mti_svvh_generic_type of Y14X10 : constant is 1;
    attribute mti_svvh_generic_type of Y14X11 : constant is 1;
    attribute mti_svvh_generic_type of Y14X12 : constant is 1;
    attribute mti_svvh_generic_type of Y14X13 : constant is 1;
    attribute mti_svvh_generic_type of Y14X14 : constant is 1;
    attribute mti_svvh_generic_type of Y14X15 : constant is 1;
    attribute mti_svvh_generic_type of Y14X16 : constant is 1;
    attribute mti_svvh_generic_type of Y14X17 : constant is 1;
    attribute mti_svvh_generic_type of Y14X18 : constant is 1;
    attribute mti_svvh_generic_type of Y14X19 : constant is 1;
    attribute mti_svvh_generic_type of Y14X20 : constant is 1;
    attribute mti_svvh_generic_type of Y14X21 : constant is 1;
    attribute mti_svvh_generic_type of Y14X22 : constant is 1;
    attribute mti_svvh_generic_type of Y14X23 : constant is 1;
    attribute mti_svvh_generic_type of Y14X24 : constant is 1;
    attribute mti_svvh_generic_type of Y14X25 : constant is 1;
    attribute mti_svvh_generic_type of Y14X26 : constant is 1;
    attribute mti_svvh_generic_type of Y14X27 : constant is 1;
    attribute mti_svvh_generic_type of Y14X28 : constant is 1;
    attribute mti_svvh_generic_type of Y15X1 : constant is 1;
    attribute mti_svvh_generic_type of Y15X2 : constant is 1;
    attribute mti_svvh_generic_type of Y15X3 : constant is 1;
    attribute mti_svvh_generic_type of Y15X4 : constant is 1;
    attribute mti_svvh_generic_type of Y15X5 : constant is 1;
    attribute mti_svvh_generic_type of Y15X6 : constant is 1;
    attribute mti_svvh_generic_type of Y15X7 : constant is 1;
    attribute mti_svvh_generic_type of Y15X8 : constant is 1;
    attribute mti_svvh_generic_type of Y15X9 : constant is 1;
    attribute mti_svvh_generic_type of Y15X10 : constant is 1;
    attribute mti_svvh_generic_type of Y15X11 : constant is 1;
    attribute mti_svvh_generic_type of Y15X12 : constant is 1;
    attribute mti_svvh_generic_type of Y15X13 : constant is 1;
    attribute mti_svvh_generic_type of Y15X14 : constant is 1;
    attribute mti_svvh_generic_type of Y15X15 : constant is 1;
    attribute mti_svvh_generic_type of Y15X16 : constant is 1;
    attribute mti_svvh_generic_type of Y15X17 : constant is 1;
    attribute mti_svvh_generic_type of Y15X18 : constant is 1;
    attribute mti_svvh_generic_type of Y15X19 : constant is 1;
    attribute mti_svvh_generic_type of Y15X20 : constant is 1;
    attribute mti_svvh_generic_type of Y15X21 : constant is 1;
    attribute mti_svvh_generic_type of Y15X22 : constant is 1;
    attribute mti_svvh_generic_type of Y15X23 : constant is 1;
    attribute mti_svvh_generic_type of Y15X24 : constant is 1;
    attribute mti_svvh_generic_type of Y15X25 : constant is 1;
    attribute mti_svvh_generic_type of Y15X26 : constant is 1;
    attribute mti_svvh_generic_type of Y15X27 : constant is 1;
    attribute mti_svvh_generic_type of Y15X28 : constant is 1;
    attribute mti_svvh_generic_type of Y16X1 : constant is 1;
    attribute mti_svvh_generic_type of Y16X2 : constant is 1;
    attribute mti_svvh_generic_type of Y16X3 : constant is 1;
    attribute mti_svvh_generic_type of Y16X4 : constant is 1;
    attribute mti_svvh_generic_type of Y16X5 : constant is 1;
    attribute mti_svvh_generic_type of Y16X6 : constant is 1;
    attribute mti_svvh_generic_type of Y16X7 : constant is 1;
    attribute mti_svvh_generic_type of Y16X8 : constant is 1;
    attribute mti_svvh_generic_type of Y16X9 : constant is 1;
    attribute mti_svvh_generic_type of Y16X10 : constant is 1;
    attribute mti_svvh_generic_type of Y16X11 : constant is 1;
    attribute mti_svvh_generic_type of Y16X12 : constant is 1;
    attribute mti_svvh_generic_type of Y16X13 : constant is 1;
    attribute mti_svvh_generic_type of Y16X14 : constant is 1;
    attribute mti_svvh_generic_type of Y16X15 : constant is 1;
    attribute mti_svvh_generic_type of Y16X16 : constant is 1;
    attribute mti_svvh_generic_type of Y16X17 : constant is 1;
    attribute mti_svvh_generic_type of Y16X18 : constant is 1;
    attribute mti_svvh_generic_type of Y16X19 : constant is 1;
    attribute mti_svvh_generic_type of Y16X20 : constant is 1;
    attribute mti_svvh_generic_type of Y16X21 : constant is 1;
    attribute mti_svvh_generic_type of Y16X22 : constant is 1;
    attribute mti_svvh_generic_type of Y16X23 : constant is 1;
    attribute mti_svvh_generic_type of Y16X24 : constant is 1;
    attribute mti_svvh_generic_type of Y16X25 : constant is 1;
    attribute mti_svvh_generic_type of Y16X26 : constant is 1;
    attribute mti_svvh_generic_type of Y16X27 : constant is 1;
    attribute mti_svvh_generic_type of Y16X28 : constant is 1;
    attribute mti_svvh_generic_type of Y17X1 : constant is 1;
    attribute mti_svvh_generic_type of Y17X2 : constant is 1;
    attribute mti_svvh_generic_type of Y17X3 : constant is 1;
    attribute mti_svvh_generic_type of Y17X4 : constant is 1;
    attribute mti_svvh_generic_type of Y17X5 : constant is 1;
    attribute mti_svvh_generic_type of Y17X6 : constant is 1;
    attribute mti_svvh_generic_type of Y17X7 : constant is 1;
    attribute mti_svvh_generic_type of Y17X8 : constant is 1;
    attribute mti_svvh_generic_type of Y17X9 : constant is 1;
    attribute mti_svvh_generic_type of Y17X10 : constant is 1;
    attribute mti_svvh_generic_type of Y17X11 : constant is 1;
    attribute mti_svvh_generic_type of Y17X12 : constant is 1;
    attribute mti_svvh_generic_type of Y17X13 : constant is 1;
    attribute mti_svvh_generic_type of Y17X14 : constant is 1;
    attribute mti_svvh_generic_type of Y17X15 : constant is 1;
    attribute mti_svvh_generic_type of Y17X16 : constant is 1;
    attribute mti_svvh_generic_type of Y17X17 : constant is 1;
    attribute mti_svvh_generic_type of Y17X18 : constant is 1;
    attribute mti_svvh_generic_type of Y17X19 : constant is 1;
    attribute mti_svvh_generic_type of Y17X20 : constant is 1;
    attribute mti_svvh_generic_type of Y17X21 : constant is 1;
    attribute mti_svvh_generic_type of Y17X22 : constant is 1;
    attribute mti_svvh_generic_type of Y17X23 : constant is 1;
    attribute mti_svvh_generic_type of Y17X24 : constant is 1;
    attribute mti_svvh_generic_type of Y17X25 : constant is 1;
    attribute mti_svvh_generic_type of Y17X26 : constant is 1;
    attribute mti_svvh_generic_type of Y17X27 : constant is 1;
    attribute mti_svvh_generic_type of Y17X28 : constant is 1;
    attribute mti_svvh_generic_type of Y18X1 : constant is 1;
    attribute mti_svvh_generic_type of Y18X2 : constant is 1;
    attribute mti_svvh_generic_type of Y18X3 : constant is 1;
    attribute mti_svvh_generic_type of Y18X4 : constant is 1;
    attribute mti_svvh_generic_type of Y18X5 : constant is 1;
    attribute mti_svvh_generic_type of Y18X6 : constant is 1;
    attribute mti_svvh_generic_type of Y18X7 : constant is 1;
    attribute mti_svvh_generic_type of Y18X8 : constant is 1;
    attribute mti_svvh_generic_type of Y18X9 : constant is 1;
    attribute mti_svvh_generic_type of Y18X10 : constant is 1;
    attribute mti_svvh_generic_type of Y18X11 : constant is 1;
    attribute mti_svvh_generic_type of Y18X12 : constant is 1;
    attribute mti_svvh_generic_type of Y18X13 : constant is 1;
    attribute mti_svvh_generic_type of Y18X14 : constant is 1;
    attribute mti_svvh_generic_type of Y18X15 : constant is 1;
    attribute mti_svvh_generic_type of Y18X16 : constant is 1;
    attribute mti_svvh_generic_type of Y18X17 : constant is 1;
    attribute mti_svvh_generic_type of Y18X18 : constant is 1;
    attribute mti_svvh_generic_type of Y18X19 : constant is 1;
    attribute mti_svvh_generic_type of Y18X20 : constant is 1;
    attribute mti_svvh_generic_type of Y18X21 : constant is 1;
    attribute mti_svvh_generic_type of Y18X22 : constant is 1;
    attribute mti_svvh_generic_type of Y18X23 : constant is 1;
    attribute mti_svvh_generic_type of Y18X24 : constant is 1;
    attribute mti_svvh_generic_type of Y18X25 : constant is 1;
    attribute mti_svvh_generic_type of Y18X26 : constant is 1;
    attribute mti_svvh_generic_type of Y18X27 : constant is 1;
    attribute mti_svvh_generic_type of Y18X28 : constant is 1;
    attribute mti_svvh_generic_type of Y19X1 : constant is 1;
    attribute mti_svvh_generic_type of Y19X2 : constant is 1;
    attribute mti_svvh_generic_type of Y19X3 : constant is 1;
    attribute mti_svvh_generic_type of Y19X4 : constant is 1;
    attribute mti_svvh_generic_type of Y19X5 : constant is 1;
    attribute mti_svvh_generic_type of Y19X6 : constant is 1;
    attribute mti_svvh_generic_type of Y19X7 : constant is 1;
    attribute mti_svvh_generic_type of Y19X8 : constant is 1;
    attribute mti_svvh_generic_type of Y19X9 : constant is 1;
    attribute mti_svvh_generic_type of Y19X10 : constant is 1;
    attribute mti_svvh_generic_type of Y19X11 : constant is 1;
    attribute mti_svvh_generic_type of Y19X12 : constant is 1;
    attribute mti_svvh_generic_type of Y19X13 : constant is 1;
    attribute mti_svvh_generic_type of Y19X14 : constant is 1;
    attribute mti_svvh_generic_type of Y19X15 : constant is 1;
    attribute mti_svvh_generic_type of Y19X16 : constant is 1;
    attribute mti_svvh_generic_type of Y19X17 : constant is 1;
    attribute mti_svvh_generic_type of Y19X18 : constant is 1;
    attribute mti_svvh_generic_type of Y19X19 : constant is 1;
    attribute mti_svvh_generic_type of Y19X20 : constant is 1;
    attribute mti_svvh_generic_type of Y19X21 : constant is 1;
    attribute mti_svvh_generic_type of Y19X22 : constant is 1;
    attribute mti_svvh_generic_type of Y19X23 : constant is 1;
    attribute mti_svvh_generic_type of Y19X24 : constant is 1;
    attribute mti_svvh_generic_type of Y19X25 : constant is 1;
    attribute mti_svvh_generic_type of Y19X26 : constant is 1;
    attribute mti_svvh_generic_type of Y19X27 : constant is 1;
    attribute mti_svvh_generic_type of Y19X28 : constant is 1;
    attribute mti_svvh_generic_type of Y20X1 : constant is 1;
    attribute mti_svvh_generic_type of Y20X2 : constant is 1;
    attribute mti_svvh_generic_type of Y20X3 : constant is 1;
    attribute mti_svvh_generic_type of Y20X4 : constant is 1;
    attribute mti_svvh_generic_type of Y20X5 : constant is 1;
    attribute mti_svvh_generic_type of Y20X6 : constant is 1;
    attribute mti_svvh_generic_type of Y20X7 : constant is 1;
    attribute mti_svvh_generic_type of Y20X8 : constant is 1;
    attribute mti_svvh_generic_type of Y20X9 : constant is 1;
    attribute mti_svvh_generic_type of Y20X10 : constant is 1;
    attribute mti_svvh_generic_type of Y20X11 : constant is 1;
    attribute mti_svvh_generic_type of Y20X12 : constant is 1;
    attribute mti_svvh_generic_type of Y20X13 : constant is 1;
    attribute mti_svvh_generic_type of Y20X14 : constant is 1;
    attribute mti_svvh_generic_type of Y20X15 : constant is 1;
    attribute mti_svvh_generic_type of Y20X16 : constant is 1;
    attribute mti_svvh_generic_type of Y20X17 : constant is 1;
    attribute mti_svvh_generic_type of Y20X18 : constant is 1;
    attribute mti_svvh_generic_type of Y20X19 : constant is 1;
    attribute mti_svvh_generic_type of Y20X20 : constant is 1;
    attribute mti_svvh_generic_type of Y20X21 : constant is 1;
    attribute mti_svvh_generic_type of Y20X22 : constant is 1;
    attribute mti_svvh_generic_type of Y20X23 : constant is 1;
    attribute mti_svvh_generic_type of Y20X24 : constant is 1;
    attribute mti_svvh_generic_type of Y20X25 : constant is 1;
    attribute mti_svvh_generic_type of Y20X26 : constant is 1;
    attribute mti_svvh_generic_type of Y20X27 : constant is 1;
    attribute mti_svvh_generic_type of Y20X28 : constant is 1;
    attribute mti_svvh_generic_type of Y21X1 : constant is 1;
    attribute mti_svvh_generic_type of Y21X2 : constant is 1;
    attribute mti_svvh_generic_type of Y21X3 : constant is 1;
    attribute mti_svvh_generic_type of Y21X4 : constant is 1;
    attribute mti_svvh_generic_type of Y21X5 : constant is 1;
    attribute mti_svvh_generic_type of Y21X6 : constant is 1;
    attribute mti_svvh_generic_type of Y21X7 : constant is 1;
    attribute mti_svvh_generic_type of Y21X8 : constant is 1;
    attribute mti_svvh_generic_type of Y21X9 : constant is 1;
    attribute mti_svvh_generic_type of Y21X10 : constant is 1;
    attribute mti_svvh_generic_type of Y21X11 : constant is 1;
    attribute mti_svvh_generic_type of Y21X12 : constant is 1;
    attribute mti_svvh_generic_type of Y21X13 : constant is 1;
    attribute mti_svvh_generic_type of Y21X14 : constant is 1;
    attribute mti_svvh_generic_type of Y21X15 : constant is 1;
    attribute mti_svvh_generic_type of Y21X16 : constant is 1;
    attribute mti_svvh_generic_type of Y21X17 : constant is 1;
    attribute mti_svvh_generic_type of Y21X18 : constant is 1;
    attribute mti_svvh_generic_type of Y21X19 : constant is 1;
    attribute mti_svvh_generic_type of Y21X20 : constant is 1;
    attribute mti_svvh_generic_type of Y21X21 : constant is 1;
    attribute mti_svvh_generic_type of Y21X22 : constant is 1;
    attribute mti_svvh_generic_type of Y21X23 : constant is 1;
    attribute mti_svvh_generic_type of Y21X24 : constant is 1;
    attribute mti_svvh_generic_type of Y21X25 : constant is 1;
    attribute mti_svvh_generic_type of Y21X26 : constant is 1;
    attribute mti_svvh_generic_type of Y21X27 : constant is 1;
    attribute mti_svvh_generic_type of Y21X28 : constant is 1;
    attribute mti_svvh_generic_type of Y22X1 : constant is 1;
    attribute mti_svvh_generic_type of Y22X2 : constant is 1;
    attribute mti_svvh_generic_type of Y22X3 : constant is 1;
    attribute mti_svvh_generic_type of Y22X4 : constant is 1;
    attribute mti_svvh_generic_type of Y22X5 : constant is 1;
    attribute mti_svvh_generic_type of Y22X6 : constant is 1;
    attribute mti_svvh_generic_type of Y22X7 : constant is 1;
    attribute mti_svvh_generic_type of Y22X8 : constant is 1;
    attribute mti_svvh_generic_type of Y22X9 : constant is 1;
    attribute mti_svvh_generic_type of Y22X10 : constant is 1;
    attribute mti_svvh_generic_type of Y22X11 : constant is 1;
    attribute mti_svvh_generic_type of Y22X12 : constant is 1;
    attribute mti_svvh_generic_type of Y22X13 : constant is 1;
    attribute mti_svvh_generic_type of Y22X14 : constant is 1;
    attribute mti_svvh_generic_type of Y22X15 : constant is 1;
    attribute mti_svvh_generic_type of Y22X16 : constant is 1;
    attribute mti_svvh_generic_type of Y22X17 : constant is 1;
    attribute mti_svvh_generic_type of Y22X18 : constant is 1;
    attribute mti_svvh_generic_type of Y22X19 : constant is 1;
    attribute mti_svvh_generic_type of Y22X20 : constant is 1;
    attribute mti_svvh_generic_type of Y22X21 : constant is 1;
    attribute mti_svvh_generic_type of Y22X22 : constant is 1;
    attribute mti_svvh_generic_type of Y22X23 : constant is 1;
    attribute mti_svvh_generic_type of Y22X24 : constant is 1;
    attribute mti_svvh_generic_type of Y22X25 : constant is 1;
    attribute mti_svvh_generic_type of Y22X26 : constant is 1;
    attribute mti_svvh_generic_type of Y22X27 : constant is 1;
    attribute mti_svvh_generic_type of Y22X28 : constant is 1;
    attribute mti_svvh_generic_type of Y23X1 : constant is 1;
    attribute mti_svvh_generic_type of Y23X2 : constant is 1;
    attribute mti_svvh_generic_type of Y23X3 : constant is 1;
    attribute mti_svvh_generic_type of Y23X4 : constant is 1;
    attribute mti_svvh_generic_type of Y23X5 : constant is 1;
    attribute mti_svvh_generic_type of Y23X6 : constant is 1;
    attribute mti_svvh_generic_type of Y23X7 : constant is 1;
    attribute mti_svvh_generic_type of Y23X8 : constant is 1;
    attribute mti_svvh_generic_type of Y23X9 : constant is 1;
    attribute mti_svvh_generic_type of Y23X10 : constant is 1;
    attribute mti_svvh_generic_type of Y23X11 : constant is 1;
    attribute mti_svvh_generic_type of Y23X12 : constant is 1;
    attribute mti_svvh_generic_type of Y23X13 : constant is 1;
    attribute mti_svvh_generic_type of Y23X14 : constant is 1;
    attribute mti_svvh_generic_type of Y23X15 : constant is 1;
    attribute mti_svvh_generic_type of Y23X16 : constant is 1;
    attribute mti_svvh_generic_type of Y23X17 : constant is 1;
    attribute mti_svvh_generic_type of Y23X18 : constant is 1;
    attribute mti_svvh_generic_type of Y23X19 : constant is 1;
    attribute mti_svvh_generic_type of Y23X20 : constant is 1;
    attribute mti_svvh_generic_type of Y23X21 : constant is 1;
    attribute mti_svvh_generic_type of Y23X22 : constant is 1;
    attribute mti_svvh_generic_type of Y23X23 : constant is 1;
    attribute mti_svvh_generic_type of Y23X24 : constant is 1;
    attribute mti_svvh_generic_type of Y23X25 : constant is 1;
    attribute mti_svvh_generic_type of Y23X26 : constant is 1;
    attribute mti_svvh_generic_type of Y23X27 : constant is 1;
    attribute mti_svvh_generic_type of Y23X28 : constant is 1;
    attribute mti_svvh_generic_type of Y24X1 : constant is 1;
    attribute mti_svvh_generic_type of Y24X2 : constant is 1;
    attribute mti_svvh_generic_type of Y24X3 : constant is 1;
    attribute mti_svvh_generic_type of Y24X4 : constant is 1;
    attribute mti_svvh_generic_type of Y24X5 : constant is 1;
    attribute mti_svvh_generic_type of Y24X6 : constant is 1;
    attribute mti_svvh_generic_type of Y24X7 : constant is 1;
    attribute mti_svvh_generic_type of Y24X8 : constant is 1;
    attribute mti_svvh_generic_type of Y24X9 : constant is 1;
    attribute mti_svvh_generic_type of Y24X10 : constant is 1;
    attribute mti_svvh_generic_type of Y24X11 : constant is 1;
    attribute mti_svvh_generic_type of Y24X12 : constant is 1;
    attribute mti_svvh_generic_type of Y24X13 : constant is 1;
    attribute mti_svvh_generic_type of Y24X14 : constant is 1;
    attribute mti_svvh_generic_type of Y24X15 : constant is 1;
    attribute mti_svvh_generic_type of Y24X16 : constant is 1;
    attribute mti_svvh_generic_type of Y24X17 : constant is 1;
    attribute mti_svvh_generic_type of Y24X18 : constant is 1;
    attribute mti_svvh_generic_type of Y24X19 : constant is 1;
    attribute mti_svvh_generic_type of Y24X20 : constant is 1;
    attribute mti_svvh_generic_type of Y24X21 : constant is 1;
    attribute mti_svvh_generic_type of Y24X22 : constant is 1;
    attribute mti_svvh_generic_type of Y24X23 : constant is 1;
    attribute mti_svvh_generic_type of Y24X24 : constant is 1;
    attribute mti_svvh_generic_type of Y24X25 : constant is 1;
    attribute mti_svvh_generic_type of Y24X26 : constant is 1;
    attribute mti_svvh_generic_type of Y24X27 : constant is 1;
    attribute mti_svvh_generic_type of Y24X28 : constant is 1;
    attribute mti_svvh_generic_type of Y25X1 : constant is 1;
    attribute mti_svvh_generic_type of Y25X2 : constant is 1;
    attribute mti_svvh_generic_type of Y25X3 : constant is 1;
    attribute mti_svvh_generic_type of Y25X4 : constant is 1;
    attribute mti_svvh_generic_type of Y25X5 : constant is 1;
    attribute mti_svvh_generic_type of Y25X6 : constant is 1;
    attribute mti_svvh_generic_type of Y25X7 : constant is 1;
    attribute mti_svvh_generic_type of Y25X8 : constant is 1;
    attribute mti_svvh_generic_type of Y25X9 : constant is 1;
    attribute mti_svvh_generic_type of Y25X10 : constant is 1;
    attribute mti_svvh_generic_type of Y25X11 : constant is 1;
    attribute mti_svvh_generic_type of Y25X12 : constant is 1;
    attribute mti_svvh_generic_type of Y25X13 : constant is 1;
    attribute mti_svvh_generic_type of Y25X14 : constant is 1;
    attribute mti_svvh_generic_type of Y25X15 : constant is 1;
    attribute mti_svvh_generic_type of Y25X16 : constant is 1;
    attribute mti_svvh_generic_type of Y25X17 : constant is 1;
    attribute mti_svvh_generic_type of Y25X18 : constant is 1;
    attribute mti_svvh_generic_type of Y25X19 : constant is 1;
    attribute mti_svvh_generic_type of Y25X20 : constant is 1;
    attribute mti_svvh_generic_type of Y25X21 : constant is 1;
    attribute mti_svvh_generic_type of Y25X22 : constant is 1;
    attribute mti_svvh_generic_type of Y25X23 : constant is 1;
    attribute mti_svvh_generic_type of Y25X24 : constant is 1;
    attribute mti_svvh_generic_type of Y25X25 : constant is 1;
    attribute mti_svvh_generic_type of Y25X26 : constant is 1;
    attribute mti_svvh_generic_type of Y25X27 : constant is 1;
    attribute mti_svvh_generic_type of Y25X28 : constant is 1;
    attribute mti_svvh_generic_type of Y26X1 : constant is 1;
    attribute mti_svvh_generic_type of Y26X2 : constant is 1;
    attribute mti_svvh_generic_type of Y26X3 : constant is 1;
    attribute mti_svvh_generic_type of Y26X4 : constant is 1;
    attribute mti_svvh_generic_type of Y26X5 : constant is 1;
    attribute mti_svvh_generic_type of Y26X6 : constant is 1;
    attribute mti_svvh_generic_type of Y26X7 : constant is 1;
    attribute mti_svvh_generic_type of Y26X8 : constant is 1;
    attribute mti_svvh_generic_type of Y26X9 : constant is 1;
    attribute mti_svvh_generic_type of Y26X10 : constant is 1;
    attribute mti_svvh_generic_type of Y26X11 : constant is 1;
    attribute mti_svvh_generic_type of Y26X12 : constant is 1;
    attribute mti_svvh_generic_type of Y26X13 : constant is 1;
    attribute mti_svvh_generic_type of Y26X14 : constant is 1;
    attribute mti_svvh_generic_type of Y26X15 : constant is 1;
    attribute mti_svvh_generic_type of Y26X16 : constant is 1;
    attribute mti_svvh_generic_type of Y26X17 : constant is 1;
    attribute mti_svvh_generic_type of Y26X18 : constant is 1;
    attribute mti_svvh_generic_type of Y26X19 : constant is 1;
    attribute mti_svvh_generic_type of Y26X20 : constant is 1;
    attribute mti_svvh_generic_type of Y26X21 : constant is 1;
    attribute mti_svvh_generic_type of Y26X22 : constant is 1;
    attribute mti_svvh_generic_type of Y26X23 : constant is 1;
    attribute mti_svvh_generic_type of Y26X24 : constant is 1;
    attribute mti_svvh_generic_type of Y26X25 : constant is 1;
    attribute mti_svvh_generic_type of Y26X26 : constant is 1;
    attribute mti_svvh_generic_type of Y26X27 : constant is 1;
    attribute mti_svvh_generic_type of Y26X28 : constant is 1;
    attribute mti_svvh_generic_type of Y27X1 : constant is 1;
    attribute mti_svvh_generic_type of Y27X2 : constant is 1;
    attribute mti_svvh_generic_type of Y27X3 : constant is 1;
    attribute mti_svvh_generic_type of Y27X4 : constant is 1;
    attribute mti_svvh_generic_type of Y27X5 : constant is 1;
    attribute mti_svvh_generic_type of Y27X6 : constant is 1;
    attribute mti_svvh_generic_type of Y27X7 : constant is 1;
    attribute mti_svvh_generic_type of Y27X8 : constant is 1;
    attribute mti_svvh_generic_type of Y27X9 : constant is 1;
    attribute mti_svvh_generic_type of Y27X10 : constant is 1;
    attribute mti_svvh_generic_type of Y27X11 : constant is 1;
    attribute mti_svvh_generic_type of Y27X12 : constant is 1;
    attribute mti_svvh_generic_type of Y27X13 : constant is 1;
    attribute mti_svvh_generic_type of Y27X14 : constant is 1;
    attribute mti_svvh_generic_type of Y27X15 : constant is 1;
    attribute mti_svvh_generic_type of Y27X16 : constant is 1;
    attribute mti_svvh_generic_type of Y27X17 : constant is 1;
    attribute mti_svvh_generic_type of Y27X18 : constant is 1;
    attribute mti_svvh_generic_type of Y27X19 : constant is 1;
    attribute mti_svvh_generic_type of Y27X20 : constant is 1;
    attribute mti_svvh_generic_type of Y27X21 : constant is 1;
    attribute mti_svvh_generic_type of Y27X22 : constant is 1;
    attribute mti_svvh_generic_type of Y27X23 : constant is 1;
    attribute mti_svvh_generic_type of Y27X24 : constant is 1;
    attribute mti_svvh_generic_type of Y27X25 : constant is 1;
    attribute mti_svvh_generic_type of Y27X26 : constant is 1;
    attribute mti_svvh_generic_type of Y27X27 : constant is 1;
    attribute mti_svvh_generic_type of Y27X28 : constant is 1;
    attribute mti_svvh_generic_type of Y28X1 : constant is 1;
    attribute mti_svvh_generic_type of Y28X2 : constant is 1;
    attribute mti_svvh_generic_type of Y28X3 : constant is 1;
    attribute mti_svvh_generic_type of Y28X4 : constant is 1;
    attribute mti_svvh_generic_type of Y28X5 : constant is 1;
    attribute mti_svvh_generic_type of Y28X6 : constant is 1;
    attribute mti_svvh_generic_type of Y28X7 : constant is 1;
    attribute mti_svvh_generic_type of Y28X8 : constant is 1;
    attribute mti_svvh_generic_type of Y28X9 : constant is 1;
    attribute mti_svvh_generic_type of Y28X10 : constant is 1;
    attribute mti_svvh_generic_type of Y28X11 : constant is 1;
    attribute mti_svvh_generic_type of Y28X12 : constant is 1;
    attribute mti_svvh_generic_type of Y28X13 : constant is 1;
    attribute mti_svvh_generic_type of Y28X14 : constant is 1;
    attribute mti_svvh_generic_type of Y28X15 : constant is 1;
    attribute mti_svvh_generic_type of Y28X16 : constant is 1;
    attribute mti_svvh_generic_type of Y28X17 : constant is 1;
    attribute mti_svvh_generic_type of Y28X18 : constant is 1;
    attribute mti_svvh_generic_type of Y28X19 : constant is 1;
    attribute mti_svvh_generic_type of Y28X20 : constant is 1;
    attribute mti_svvh_generic_type of Y28X21 : constant is 1;
    attribute mti_svvh_generic_type of Y28X22 : constant is 1;
    attribute mti_svvh_generic_type of Y28X23 : constant is 1;
    attribute mti_svvh_generic_type of Y28X24 : constant is 1;
    attribute mti_svvh_generic_type of Y28X25 : constant is 1;
    attribute mti_svvh_generic_type of Y28X26 : constant is 1;
    attribute mti_svvh_generic_type of Y28X27 : constant is 1;
    attribute mti_svvh_generic_type of Y28X28 : constant is 1;
    attribute mti_svvh_generic_type of Y29X1 : constant is 1;
    attribute mti_svvh_generic_type of Y29X2 : constant is 1;
    attribute mti_svvh_generic_type of Y29X3 : constant is 1;
    attribute mti_svvh_generic_type of Y29X4 : constant is 1;
    attribute mti_svvh_generic_type of Y29X5 : constant is 1;
    attribute mti_svvh_generic_type of Y29X6 : constant is 1;
    attribute mti_svvh_generic_type of Y29X7 : constant is 1;
    attribute mti_svvh_generic_type of Y29X8 : constant is 1;
    attribute mti_svvh_generic_type of Y29X9 : constant is 1;
    attribute mti_svvh_generic_type of Y29X10 : constant is 1;
    attribute mti_svvh_generic_type of Y29X11 : constant is 1;
    attribute mti_svvh_generic_type of Y29X12 : constant is 1;
    attribute mti_svvh_generic_type of Y29X13 : constant is 1;
    attribute mti_svvh_generic_type of Y29X14 : constant is 1;
    attribute mti_svvh_generic_type of Y29X15 : constant is 1;
    attribute mti_svvh_generic_type of Y29X16 : constant is 1;
    attribute mti_svvh_generic_type of Y29X17 : constant is 1;
    attribute mti_svvh_generic_type of Y29X18 : constant is 1;
    attribute mti_svvh_generic_type of Y29X19 : constant is 1;
    attribute mti_svvh_generic_type of Y29X20 : constant is 1;
    attribute mti_svvh_generic_type of Y29X21 : constant is 1;
    attribute mti_svvh_generic_type of Y29X22 : constant is 1;
    attribute mti_svvh_generic_type of Y29X23 : constant is 1;
    attribute mti_svvh_generic_type of Y29X24 : constant is 1;
    attribute mti_svvh_generic_type of Y29X25 : constant is 1;
    attribute mti_svvh_generic_type of Y29X26 : constant is 1;
    attribute mti_svvh_generic_type of Y29X27 : constant is 1;
    attribute mti_svvh_generic_type of Y29X28 : constant is 1;
    attribute mti_svvh_generic_type of Y30X1 : constant is 1;
    attribute mti_svvh_generic_type of Y30X2 : constant is 1;
    attribute mti_svvh_generic_type of Y30X3 : constant is 1;
    attribute mti_svvh_generic_type of Y30X4 : constant is 1;
    attribute mti_svvh_generic_type of Y30X5 : constant is 1;
    attribute mti_svvh_generic_type of Y30X6 : constant is 1;
    attribute mti_svvh_generic_type of Y30X7 : constant is 1;
    attribute mti_svvh_generic_type of Y30X8 : constant is 1;
    attribute mti_svvh_generic_type of Y30X9 : constant is 1;
    attribute mti_svvh_generic_type of Y30X10 : constant is 1;
    attribute mti_svvh_generic_type of Y30X11 : constant is 1;
    attribute mti_svvh_generic_type of Y30X12 : constant is 1;
    attribute mti_svvh_generic_type of Y30X13 : constant is 1;
    attribute mti_svvh_generic_type of Y30X14 : constant is 1;
    attribute mti_svvh_generic_type of Y30X15 : constant is 1;
    attribute mti_svvh_generic_type of Y30X16 : constant is 1;
    attribute mti_svvh_generic_type of Y30X17 : constant is 1;
    attribute mti_svvh_generic_type of Y30X18 : constant is 1;
    attribute mti_svvh_generic_type of Y30X19 : constant is 1;
    attribute mti_svvh_generic_type of Y30X20 : constant is 1;
    attribute mti_svvh_generic_type of Y30X21 : constant is 1;
    attribute mti_svvh_generic_type of Y30X22 : constant is 1;
    attribute mti_svvh_generic_type of Y30X23 : constant is 1;
    attribute mti_svvh_generic_type of Y30X24 : constant is 1;
    attribute mti_svvh_generic_type of Y30X25 : constant is 1;
    attribute mti_svvh_generic_type of Y30X26 : constant is 1;
    attribute mti_svvh_generic_type of Y30X27 : constant is 1;
    attribute mti_svvh_generic_type of Y30X28 : constant is 1;
    attribute mti_svvh_generic_type of Y31X1 : constant is 1;
    attribute mti_svvh_generic_type of Y31X2 : constant is 1;
    attribute mti_svvh_generic_type of Y31X3 : constant is 1;
    attribute mti_svvh_generic_type of Y31X4 : constant is 1;
    attribute mti_svvh_generic_type of Y31X5 : constant is 1;
    attribute mti_svvh_generic_type of Y31X6 : constant is 1;
    attribute mti_svvh_generic_type of Y31X7 : constant is 1;
    attribute mti_svvh_generic_type of Y31X8 : constant is 1;
    attribute mti_svvh_generic_type of Y31X9 : constant is 1;
    attribute mti_svvh_generic_type of Y31X10 : constant is 1;
    attribute mti_svvh_generic_type of Y31X11 : constant is 1;
    attribute mti_svvh_generic_type of Y31X12 : constant is 1;
    attribute mti_svvh_generic_type of Y31X13 : constant is 1;
    attribute mti_svvh_generic_type of Y31X14 : constant is 1;
    attribute mti_svvh_generic_type of Y31X15 : constant is 1;
    attribute mti_svvh_generic_type of Y31X16 : constant is 1;
    attribute mti_svvh_generic_type of Y31X17 : constant is 1;
    attribute mti_svvh_generic_type of Y31X18 : constant is 1;
    attribute mti_svvh_generic_type of Y31X19 : constant is 1;
    attribute mti_svvh_generic_type of Y31X20 : constant is 1;
    attribute mti_svvh_generic_type of Y31X21 : constant is 1;
    attribute mti_svvh_generic_type of Y31X22 : constant is 1;
    attribute mti_svvh_generic_type of Y31X23 : constant is 1;
    attribute mti_svvh_generic_type of Y31X24 : constant is 1;
    attribute mti_svvh_generic_type of Y31X25 : constant is 1;
    attribute mti_svvh_generic_type of Y31X26 : constant is 1;
    attribute mti_svvh_generic_type of Y31X27 : constant is 1;
    attribute mti_svvh_generic_type of Y31X28 : constant is 1;
    attribute mti_svvh_generic_type of Y32X1 : constant is 1;
    attribute mti_svvh_generic_type of Y32X2 : constant is 1;
    attribute mti_svvh_generic_type of Y32X3 : constant is 1;
    attribute mti_svvh_generic_type of Y32X4 : constant is 1;
    attribute mti_svvh_generic_type of Y32X5 : constant is 1;
    attribute mti_svvh_generic_type of Y32X6 : constant is 1;
    attribute mti_svvh_generic_type of Y32X7 : constant is 1;
    attribute mti_svvh_generic_type of Y32X8 : constant is 1;
    attribute mti_svvh_generic_type of Y32X9 : constant is 1;
    attribute mti_svvh_generic_type of Y32X10 : constant is 1;
    attribute mti_svvh_generic_type of Y32X11 : constant is 1;
    attribute mti_svvh_generic_type of Y32X12 : constant is 1;
    attribute mti_svvh_generic_type of Y32X13 : constant is 1;
    attribute mti_svvh_generic_type of Y32X14 : constant is 1;
    attribute mti_svvh_generic_type of Y32X15 : constant is 1;
    attribute mti_svvh_generic_type of Y32X16 : constant is 1;
    attribute mti_svvh_generic_type of Y32X17 : constant is 1;
    attribute mti_svvh_generic_type of Y32X18 : constant is 1;
    attribute mti_svvh_generic_type of Y32X19 : constant is 1;
    attribute mti_svvh_generic_type of Y32X20 : constant is 1;
    attribute mti_svvh_generic_type of Y32X21 : constant is 1;
    attribute mti_svvh_generic_type of Y32X22 : constant is 1;
    attribute mti_svvh_generic_type of Y32X23 : constant is 1;
    attribute mti_svvh_generic_type of Y32X24 : constant is 1;
    attribute mti_svvh_generic_type of Y32X25 : constant is 1;
    attribute mti_svvh_generic_type of Y32X26 : constant is 1;
    attribute mti_svvh_generic_type of Y32X27 : constant is 1;
    attribute mti_svvh_generic_type of Y32X28 : constant is 1;
    attribute mti_svvh_generic_type of Y33X1 : constant is 1;
    attribute mti_svvh_generic_type of Y33X2 : constant is 1;
    attribute mti_svvh_generic_type of Y33X3 : constant is 1;
    attribute mti_svvh_generic_type of Y33X4 : constant is 1;
    attribute mti_svvh_generic_type of Y33X5 : constant is 1;
    attribute mti_svvh_generic_type of Y33X6 : constant is 1;
    attribute mti_svvh_generic_type of Y33X7 : constant is 1;
    attribute mti_svvh_generic_type of Y33X8 : constant is 1;
    attribute mti_svvh_generic_type of Y33X9 : constant is 1;
    attribute mti_svvh_generic_type of Y33X10 : constant is 1;
    attribute mti_svvh_generic_type of Y33X11 : constant is 1;
    attribute mti_svvh_generic_type of Y33X12 : constant is 1;
    attribute mti_svvh_generic_type of Y33X13 : constant is 1;
    attribute mti_svvh_generic_type of Y33X14 : constant is 1;
    attribute mti_svvh_generic_type of Y33X15 : constant is 1;
    attribute mti_svvh_generic_type of Y33X16 : constant is 1;
    attribute mti_svvh_generic_type of Y33X17 : constant is 1;
    attribute mti_svvh_generic_type of Y33X18 : constant is 1;
    attribute mti_svvh_generic_type of Y33X19 : constant is 1;
    attribute mti_svvh_generic_type of Y33X20 : constant is 1;
    attribute mti_svvh_generic_type of Y33X21 : constant is 1;
    attribute mti_svvh_generic_type of Y33X22 : constant is 1;
    attribute mti_svvh_generic_type of Y33X23 : constant is 1;
    attribute mti_svvh_generic_type of Y33X24 : constant is 1;
    attribute mti_svvh_generic_type of Y33X25 : constant is 1;
    attribute mti_svvh_generic_type of Y33X26 : constant is 1;
    attribute mti_svvh_generic_type of Y33X27 : constant is 1;
    attribute mti_svvh_generic_type of Y33X28 : constant is 1;
    attribute mti_svvh_generic_type of Y34X1 : constant is 1;
    attribute mti_svvh_generic_type of Y34X2 : constant is 1;
    attribute mti_svvh_generic_type of Y34X3 : constant is 1;
    attribute mti_svvh_generic_type of Y34X4 : constant is 1;
    attribute mti_svvh_generic_type of Y34X5 : constant is 1;
    attribute mti_svvh_generic_type of Y34X6 : constant is 1;
    attribute mti_svvh_generic_type of Y34X7 : constant is 1;
    attribute mti_svvh_generic_type of Y34X8 : constant is 1;
    attribute mti_svvh_generic_type of Y34X9 : constant is 1;
    attribute mti_svvh_generic_type of Y34X10 : constant is 1;
    attribute mti_svvh_generic_type of Y34X11 : constant is 1;
    attribute mti_svvh_generic_type of Y34X12 : constant is 1;
    attribute mti_svvh_generic_type of Y34X13 : constant is 1;
    attribute mti_svvh_generic_type of Y34X14 : constant is 1;
    attribute mti_svvh_generic_type of Y34X15 : constant is 1;
    attribute mti_svvh_generic_type of Y34X16 : constant is 1;
    attribute mti_svvh_generic_type of Y34X17 : constant is 1;
    attribute mti_svvh_generic_type of Y34X18 : constant is 1;
    attribute mti_svvh_generic_type of Y34X19 : constant is 1;
    attribute mti_svvh_generic_type of Y34X20 : constant is 1;
    attribute mti_svvh_generic_type of Y34X21 : constant is 1;
    attribute mti_svvh_generic_type of Y34X22 : constant is 1;
    attribute mti_svvh_generic_type of Y34X23 : constant is 1;
    attribute mti_svvh_generic_type of Y34X24 : constant is 1;
    attribute mti_svvh_generic_type of Y34X25 : constant is 1;
    attribute mti_svvh_generic_type of Y34X26 : constant is 1;
    attribute mti_svvh_generic_type of Y34X27 : constant is 1;
    attribute mti_svvh_generic_type of Y34X28 : constant is 1;
    attribute mti_svvh_generic_type of Y35X1 : constant is 1;
    attribute mti_svvh_generic_type of Y35X2 : constant is 1;
    attribute mti_svvh_generic_type of Y35X3 : constant is 1;
    attribute mti_svvh_generic_type of Y35X4 : constant is 1;
    attribute mti_svvh_generic_type of Y35X5 : constant is 1;
    attribute mti_svvh_generic_type of Y35X6 : constant is 1;
    attribute mti_svvh_generic_type of Y35X7 : constant is 1;
    attribute mti_svvh_generic_type of Y35X8 : constant is 1;
    attribute mti_svvh_generic_type of Y35X9 : constant is 1;
    attribute mti_svvh_generic_type of Y35X10 : constant is 1;
    attribute mti_svvh_generic_type of Y35X11 : constant is 1;
    attribute mti_svvh_generic_type of Y35X12 : constant is 1;
    attribute mti_svvh_generic_type of Y35X13 : constant is 1;
    attribute mti_svvh_generic_type of Y35X14 : constant is 1;
    attribute mti_svvh_generic_type of Y35X15 : constant is 1;
    attribute mti_svvh_generic_type of Y35X16 : constant is 1;
    attribute mti_svvh_generic_type of Y35X17 : constant is 1;
    attribute mti_svvh_generic_type of Y35X18 : constant is 1;
    attribute mti_svvh_generic_type of Y35X19 : constant is 1;
    attribute mti_svvh_generic_type of Y35X20 : constant is 1;
    attribute mti_svvh_generic_type of Y35X21 : constant is 1;
    attribute mti_svvh_generic_type of Y35X22 : constant is 1;
    attribute mti_svvh_generic_type of Y35X23 : constant is 1;
    attribute mti_svvh_generic_type of Y35X24 : constant is 1;
    attribute mti_svvh_generic_type of Y35X25 : constant is 1;
    attribute mti_svvh_generic_type of Y35X26 : constant is 1;
    attribute mti_svvh_generic_type of Y35X27 : constant is 1;
    attribute mti_svvh_generic_type of Y35X28 : constant is 1;
    attribute mti_svvh_generic_type of YY0XX0 : constant is 1;
    attribute mti_svvh_generic_type of YY0XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY0XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY0XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY0XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY0XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY0XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY0XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY0XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY0XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY0XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY0XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY0XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY0XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY0XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY0XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY0XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY0XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY0XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY0XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY0XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY0XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY0XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY0XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY0XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY0XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY0XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY0XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY0XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY1XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY1XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY1XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY1XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY1XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY1XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY1XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY1XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY1XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY1XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY1XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY1XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY1XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY1XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY1XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY1XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY1XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY1XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY1XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY1XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY1XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY1XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY1XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY1XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY1XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY1XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY1XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY1XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY2XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY2XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY2XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY2XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY2XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY2XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY2XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY2XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY2XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY2XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY2XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY2XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY2XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY2XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY2XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY2XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY2XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY2XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY2XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY2XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY2XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY2XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY2XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY2XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY2XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY2XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY2XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY2XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY3XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY3XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY3XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY3XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY3XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY3XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY3XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY3XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY3XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY3XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY3XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY3XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY3XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY3XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY3XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY3XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY3XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY3XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY3XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY3XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY3XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY3XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY3XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY3XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY3XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY3XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY3XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY3XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY4XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY4XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY4XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY4XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY4XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY4XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY4XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY4XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY4XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY4XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY4XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY4XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY4XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY4XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY4XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY4XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY4XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY4XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY4XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY4XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY4XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY4XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY4XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY4XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY4XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY4XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY4XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY4XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY5XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY5XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY5XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY5XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY5XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY5XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY5XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY5XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY5XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY5XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY5XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY5XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY5XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY5XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY5XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY5XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY5XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY5XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY5XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY5XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY5XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY5XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY5XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY5XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY5XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY5XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY5XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY5XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY6XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY6XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY6XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY6XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY6XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY6XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY6XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY6XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY6XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY6XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY6XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY6XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY6XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY6XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY6XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY6XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY6XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY6XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY6XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY6XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY6XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY6XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY6XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY6XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY6XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY6XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY6XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY6XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY7XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY7XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY7XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY7XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY7XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY7XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY7XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY7XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY7XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY7XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY7XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY7XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY7XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY7XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY7XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY7XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY7XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY7XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY7XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY7XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY7XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY7XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY7XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY7XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY7XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY7XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY7XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY7XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY8XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY8XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY8XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY8XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY8XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY8XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY8XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY8XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY8XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY8XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY8XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY8XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY8XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY8XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY8XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY8XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY8XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY8XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY8XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY8XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY8XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY8XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY8XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY8XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY8XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY8XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY8XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY8XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY9XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY9XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY9XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY9XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY9XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY9XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY9XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY9XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY9XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY9XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY9XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY9XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY9XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY9XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY9XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY9XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY9XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY9XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY9XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY9XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY9XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY9XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY9XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY9XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY9XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY9XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY9XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY9XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY10XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY10XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY10XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY10XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY10XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY10XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY10XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY10XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY10XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY10XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY10XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY10XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY10XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY10XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY10XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY10XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY10XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY10XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY10XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY10XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY10XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY10XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY10XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY10XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY10XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY10XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY10XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY10XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY11XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY11XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY11XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY11XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY11XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY11XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY11XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY11XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY11XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY11XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY11XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY11XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY11XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY11XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY11XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY11XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY11XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY11XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY11XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY11XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY11XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY11XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY11XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY11XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY11XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY11XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY11XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY11XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY12XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY12XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY12XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY12XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY12XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY12XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY12XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY12XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY12XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY12XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY12XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY12XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY12XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY12XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY12XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY12XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY12XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY12XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY12XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY12XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY12XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY12XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY12XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY12XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY12XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY12XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY12XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY12XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY13XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY13XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY13XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY13XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY13XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY13XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY13XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY13XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY13XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY13XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY13XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY13XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY13XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY13XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY13XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY13XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY13XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY13XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY13XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY13XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY13XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY13XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY13XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY13XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY13XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY13XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY13XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY13XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY14XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY14XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY14XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY14XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY14XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY14XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY14XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY14XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY14XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY14XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY14XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY14XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY14XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY14XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY14XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY14XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY14XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY14XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY14XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY14XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY14XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY14XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY14XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY14XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY14XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY14XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY14XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY14XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY15XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY15XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY15XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY15XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY15XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY15XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY15XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY15XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY15XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY15XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY15XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY15XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY15XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY15XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY15XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY15XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY15XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY15XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY15XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY15XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY15XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY15XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY15XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY15XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY15XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY15XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY15XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY15XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY16XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY16XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY16XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY16XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY16XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY16XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY16XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY16XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY16XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY16XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY16XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY16XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY16XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY16XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY16XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY16XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY16XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY16XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY16XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY16XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY16XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY16XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY16XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY16XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY16XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY16XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY16XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY16XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY17XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY17XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY17XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY17XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY17XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY17XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY17XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY17XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY17XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY17XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY17XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY17XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY17XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY17XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY17XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY17XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY17XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY17XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY17XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY17XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY17XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY17XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY17XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY17XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY17XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY17XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY17XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY17XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY18XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY18XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY18XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY18XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY18XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY18XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY18XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY18XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY18XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY18XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY18XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY18XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY18XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY18XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY18XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY18XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY18XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY18XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY18XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY18XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY18XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY18XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY18XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY18XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY18XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY18XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY18XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY18XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY19XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY19XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY19XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY19XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY19XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY19XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY19XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY19XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY19XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY19XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY19XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY19XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY19XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY19XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY19XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY19XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY19XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY19XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY19XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY19XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY19XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY19XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY19XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY19XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY19XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY19XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY19XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY19XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY20XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY20XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY20XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY20XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY20XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY20XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY20XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY20XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY20XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY20XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY20XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY20XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY20XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY20XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY20XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY20XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY20XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY20XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY20XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY20XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY20XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY20XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY20XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY20XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY20XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY20XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY20XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY20XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY21XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY21XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY21XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY21XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY21XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY21XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY21XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY21XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY21XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY21XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY21XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY21XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY21XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY21XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY21XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY21XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY21XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY21XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY21XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY21XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY21XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY21XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY21XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY21XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY21XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY21XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY21XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY21XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY22XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY22XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY22XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY22XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY22XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY22XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY22XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY22XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY22XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY22XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY22XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY22XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY22XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY22XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY22XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY22XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY22XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY22XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY22XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY22XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY22XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY22XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY22XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY22XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY22XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY22XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY22XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY22XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY23XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY23XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY23XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY23XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY23XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY23XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY23XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY23XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY23XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY23XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY23XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY23XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY23XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY23XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY23XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY23XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY23XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY23XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY23XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY23XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY23XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY23XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY23XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY23XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY23XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY23XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY23XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY23XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY24XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY24XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY24XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY24XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY24XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY24XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY24XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY24XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY24XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY24XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY24XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY24XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY24XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY24XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY24XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY24XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY24XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY24XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY24XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY24XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY24XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY24XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY24XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY24XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY24XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY24XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY24XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY24XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY25XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY25XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY25XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY25XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY25XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY25XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY25XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY25XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY25XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY25XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY25XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY25XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY25XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY25XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY25XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY25XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY25XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY25XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY25XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY25XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY25XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY25XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY25XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY25XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY25XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY25XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY25XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY25XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY26XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY26XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY26XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY26XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY26XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY26XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY26XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY26XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY26XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY26XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY26XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY26XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY26XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY26XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY26XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY26XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY26XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY26XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY26XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY26XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY26XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY26XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY26XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY26XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY26XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY26XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY26XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY26XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY27XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY27XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY27XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY27XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY27XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY27XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY27XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY27XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY27XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY27XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY27XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY27XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY27XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY27XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY27XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY27XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY27XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY27XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY27XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY27XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY27XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY27XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY27XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY27XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY27XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY27XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY27XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY27XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY28XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY28XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY28XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY28XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY28XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY28XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY28XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY28XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY28XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY28XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY28XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY28XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY28XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY28XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY28XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY28XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY28XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY28XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY28XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY28XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY28XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY28XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY28XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY28XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY28XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY28XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY28XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY28XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY29XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY29XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY29XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY29XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY29XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY29XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY29XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY29XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY29XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY29XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY29XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY29XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY29XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY29XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY29XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY29XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY29XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY29XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY29XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY29XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY29XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY29XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY29XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY29XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY29XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY29XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY29XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY29XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY30XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY30XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY30XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY30XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY30XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY30XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY30XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY30XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY30XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY30XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY30XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY30XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY30XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY30XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY30XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY30XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY30XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY30XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY30XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY30XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY30XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY30XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY30XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY30XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY30XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY30XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY30XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY30XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY31XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY31XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY31XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY31XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY31XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY31XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY31XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY31XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY31XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY31XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY31XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY31XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY31XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY31XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY31XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY31XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY31XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY31XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY31XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY31XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY31XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY31XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY31XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY31XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY31XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY31XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY31XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY31XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY32XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY32XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY32XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY32XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY32XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY32XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY32XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY32XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY32XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY32XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY32XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY32XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY32XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY32XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY32XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY32XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY32XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY32XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY32XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY32XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY32XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY32XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY32XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY32XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY32XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY32XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY32XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY32XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY33XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY33XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY33XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY33XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY33XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY33XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY33XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY33XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY33XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY33XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY33XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY33XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY33XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY33XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY33XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY33XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY33XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY33XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY33XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY33XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY33XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY33XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY33XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY33XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY33XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY33XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY33XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY33XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY34XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY34XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY34XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY34XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY34XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY34XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY34XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY34XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY34XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY34XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY34XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY34XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY34XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY34XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY34XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY34XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY34XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY34XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY34XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY34XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY34XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY34XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY34XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY34XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY34XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY34XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY34XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY34XX28 : constant is 1;
    attribute mti_svvh_generic_type of YY35XX1 : constant is 1;
    attribute mti_svvh_generic_type of YY35XX2 : constant is 1;
    attribute mti_svvh_generic_type of YY35XX3 : constant is 1;
    attribute mti_svvh_generic_type of YY35XX4 : constant is 1;
    attribute mti_svvh_generic_type of YY35XX5 : constant is 1;
    attribute mti_svvh_generic_type of YY35XX6 : constant is 1;
    attribute mti_svvh_generic_type of YY35XX7 : constant is 1;
    attribute mti_svvh_generic_type of YY35XX8 : constant is 1;
    attribute mti_svvh_generic_type of YY35XX9 : constant is 1;
    attribute mti_svvh_generic_type of YY35XX10 : constant is 1;
    attribute mti_svvh_generic_type of YY35XX11 : constant is 1;
    attribute mti_svvh_generic_type of YY35XX12 : constant is 1;
    attribute mti_svvh_generic_type of YY35XX13 : constant is 1;
    attribute mti_svvh_generic_type of YY35XX14 : constant is 1;
    attribute mti_svvh_generic_type of YY35XX15 : constant is 1;
    attribute mti_svvh_generic_type of YY35XX16 : constant is 1;
    attribute mti_svvh_generic_type of YY35XX17 : constant is 1;
    attribute mti_svvh_generic_type of YY35XX18 : constant is 1;
    attribute mti_svvh_generic_type of YY35XX19 : constant is 1;
    attribute mti_svvh_generic_type of YY35XX20 : constant is 1;
    attribute mti_svvh_generic_type of YY35XX21 : constant is 1;
    attribute mti_svvh_generic_type of YY35XX22 : constant is 1;
    attribute mti_svvh_generic_type of YY35XX23 : constant is 1;
    attribute mti_svvh_generic_type of YY35XX24 : constant is 1;
    attribute mti_svvh_generic_type of YY35XX25 : constant is 1;
    attribute mti_svvh_generic_type of YY35XX26 : constant is 1;
    attribute mti_svvh_generic_type of YY35XX27 : constant is 1;
    attribute mti_svvh_generic_type of YY35XX28 : constant is 1;
end FFXII_LB_Cursor;
