library verilog;
use verilog.vl_types.all;
entity ksa_vlg_vec_tst is
end ksa_vlg_vec_tst;
