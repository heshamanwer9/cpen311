// DE2_QSYS.v

// Generated using ACDS version 13.0sp1 232 at 2017.04.04.15:33:00

`timescale 1 ps / 1 ps
module DE2_QSYS (
		output wire [31:0] audio2fifo_0_data_divfrec_export,                  //                  audio2fifo_0_data_divfrec.export
		input  wire        audio2fifo_0_empty_export,                         //                         audio2fifo_0_empty.export
		input  wire        audio2fifo_0_fifo_full_export,                     //                     audio2fifo_0_fifo_full.export
		input  wire [11:0] audio2fifo_0_fifo_used_export,                     //                     audio2fifo_0_fifo_used.export
		output wire [31:0] audio2fifo_0_out_data_audio_export,                //                audio2fifo_0_out_data_audio.export
		output wire        audio2fifo_0_out_pause_export,                     //                     audio2fifo_0_out_pause.export
		output wire        audio2fifo_0_out_stop_export,                      //                      audio2fifo_0_out_stop.export
		output wire        audio2fifo_0_wrclk_export,                         //                         audio2fifo_0_wrclk.export
		output wire        audio2fifo_0_wrreq_export,                         //                         audio2fifo_0_wrreq.export
		output wire        audio_sel_export,                                  //                                  audio_sel.export
		input  wire        clk_clk,                                           //                                        clk.clk
		output wire [31:0] div_freq_export,                                   //                                   div_freq.export
		input  wire [3:0]  key_external_connection_export,                    //                    key_external_connection.export
		input  wire [31:0] keyboard_keys_export,                              //                              keyboard_keys.export
		output wire [3:0]  modulation_selector_export,                        //                        modulation_selector.export
		input  wire [31:0] mouse_pos_export,                                  //                                  mouse_pos.export
		input  wire        reset_reset_n,                                     //                                      reset.reset_n
		output wire [11:0] sdram_wire_addr,                                   //                                 sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                                     //                                           .ba
		output wire        sdram_wire_cas_n,                                  //                                           .cas_n
		output wire        sdram_wire_cke,                                    //                                           .cke
		output wire        sdram_wire_cs_n,                                   //                                           .cs_n
		inout  wire [15:0] sdram_wire_dq,                                     //                                           .dq
		output wire [1:0]  sdram_wire_dqm,                                    //                                           .dqm
		output wire        sdram_wire_ras_n,                                  //                                           .ras_n
		output wire        sdram_wire_we_n,                                   //                                           .we_n
		output wire [7:0]  signal_selector_export,                            //                            signal_selector.export
		input  wire        vga_alt_vip_itc_0_clocked_video_vid_clk,           //            vga_alt_vip_itc_0_clocked_video.vid_clk
		output wire [23:0] vga_alt_vip_itc_0_clocked_video_vid_data,          //                                           .vid_data
		output wire        vga_alt_vip_itc_0_clocked_video_underflow,         //                                           .underflow
		output wire        vga_alt_vip_itc_0_clocked_video_vid_datavalid,     //                                           .vid_datavalid
		output wire        vga_alt_vip_itc_0_clocked_video_vid_v_sync,        //                                           .vid_v_sync
		output wire        vga_alt_vip_itc_0_clocked_video_vid_h_sync,        //                                           .vid_h_sync
		output wire        vga_alt_vip_itc_0_clocked_video_vid_f,             //                                           .vid_f
		output wire        vga_alt_vip_itc_0_clocked_video_vid_h,             //                                           .vid_h
		output wire        vga_alt_vip_itc_0_clocked_video_vid_v,             //                                           .vid_v
		output wire        vga_vga_clk_clk,                                   //                                vga_vga_clk.clk
		input  wire        clk_25_in_clk,                                     //                                  clk_25_in.clk
		input  wire        clk_40_in_clk,                                     //                                  clk_40_in.clk
		input  wire        cpu_clk_for_sdram_clk,                             //                          cpu_clk_for_sdram.clk
		input  wire        lfsr_clk_interrupt_gen_external_connection_export, // lfsr_clk_interrupt_gen_external_connection.export
		input  wire [31:0] lfsr_val_external_connection_export,               //               lfsr_val_external_connection.export
		output wire [31:0] dds_increment_external_connection_export           //          dds_increment_external_connection.export
	);

	wire          cpu_data_master_waitrequest;                                                                      // cpu_data_master_translator:av_waitrequest -> cpu:d_waitrequest
	wire   [31:0] cpu_data_master_writedata;                                                                        // cpu:d_writedata -> cpu_data_master_translator:av_writedata
	wire   [24:0] cpu_data_master_address;                                                                          // cpu:d_address -> cpu_data_master_translator:av_address
	wire          cpu_data_master_write;                                                                            // cpu:d_write -> cpu_data_master_translator:av_write
	wire          cpu_data_master_read;                                                                             // cpu:d_read -> cpu_data_master_translator:av_read
	wire   [31:0] cpu_data_master_readdata;                                                                         // cpu_data_master_translator:av_readdata -> cpu:d_readdata
	wire          cpu_data_master_debugaccess;                                                                      // cpu:jtag_debug_module_debugaccess_to_roms -> cpu_data_master_translator:av_debugaccess
	wire    [3:0] cpu_data_master_byteenable;                                                                       // cpu:d_byteenable -> cpu_data_master_translator:av_byteenable
	wire          vga_to_sdram_waitrequest;                                                                         // vga_to_sdram_translator:av_waitrequest -> vga:to_sdram_waitrequest
	wire    [5:0] vga_to_sdram_burstcount;                                                                          // vga:to_sdram_burstcount -> vga_to_sdram_translator:av_burstcount
	wire   [31:0] vga_to_sdram_address;                                                                             // vga:to_sdram_address -> vga_to_sdram_translator:av_address
	wire          vga_to_sdram_read;                                                                                // vga:to_sdram_read -> vga_to_sdram_translator:av_read
	wire   [31:0] vga_to_sdram_readdata;                                                                            // vga_to_sdram_translator:av_readdata -> vga:to_sdram_readdata
	wire          vga_to_sdram_readdatavalid;                                                                       // vga_to_sdram_translator:av_readdatavalid -> vga:to_sdram_readdatavalid
	wire          cpu_instruction_master_waitrequest;                                                               // cpu_instruction_master_translator:av_waitrequest -> cpu:i_waitrequest
	wire   [24:0] cpu_instruction_master_address;                                                                   // cpu:i_address -> cpu_instruction_master_translator:av_address
	wire          cpu_instruction_master_read;                                                                      // cpu:i_read -> cpu_instruction_master_translator:av_read
	wire   [31:0] cpu_instruction_master_readdata;                                                                  // cpu_instruction_master_translator:av_readdata -> cpu:i_readdata
	wire          cpu_instruction_master_readdatavalid;                                                             // cpu_instruction_master_translator:av_readdatavalid -> cpu:i_readdatavalid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                           // jtag_uart:av_waitrequest -> jtag_uart_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                             // jtag_uart_avalon_jtag_slave_translator:av_writedata -> jtag_uart:av_writedata
	wire    [0:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                               // jtag_uart_avalon_jtag_slave_translator:av_address -> jtag_uart:av_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                            // jtag_uart_avalon_jtag_slave_translator:av_chipselect -> jtag_uart:av_chipselect
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                 // jtag_uart_avalon_jtag_slave_translator:av_write -> jtag_uart:av_write_n
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                  // jtag_uart_avalon_jtag_slave_translator:av_read -> jtag_uart:av_read_n
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                              // jtag_uart:av_readdata -> jtag_uart_avalon_jtag_slave_translator:av_readdata
	wire    [0:0] sysid_qsys_control_slave_translator_avalon_anti_slave_0_address;                                  // sysid_qsys_control_slave_translator:av_address -> sysid_qsys:address
	wire   [31:0] sysid_qsys_control_slave_translator_avalon_anti_slave_0_readdata;                                 // sysid_qsys:readdata -> sysid_qsys_control_slave_translator:av_readdata
	wire   [31:0] audio_data_fregen_s1_translator_avalon_anti_slave_0_writedata;                                    // audio_data_fregen_s1_translator:av_writedata -> audio:data_fregen_s1_writedata
	wire    [1:0] audio_data_fregen_s1_translator_avalon_anti_slave_0_address;                                      // audio_data_fregen_s1_translator:av_address -> audio:data_fregen_s1_address
	wire          audio_data_fregen_s1_translator_avalon_anti_slave_0_chipselect;                                   // audio_data_fregen_s1_translator:av_chipselect -> audio:data_fregen_s1_chipselect
	wire          audio_data_fregen_s1_translator_avalon_anti_slave_0_write;                                        // audio_data_fregen_s1_translator:av_write -> audio:data_fregen_s1_write_n
	wire   [31:0] audio_data_fregen_s1_translator_avalon_anti_slave_0_readdata;                                     // audio:data_fregen_s1_readdata -> audio_data_fregen_s1_translator:av_readdata
	wire    [1:0] audio_empty_s1_translator_avalon_anti_slave_0_address;                                            // audio_empty_s1_translator:av_address -> audio:empty_s1_address
	wire   [31:0] audio_empty_s1_translator_avalon_anti_slave_0_readdata;                                           // audio:empty_s1_readdata -> audio_empty_s1_translator:av_readdata
	wire    [1:0] audio_fifo_full_s1_translator_avalon_anti_slave_0_address;                                        // audio_fifo_full_s1_translator:av_address -> audio:fifo_full_s1_address
	wire   [31:0] audio_fifo_full_s1_translator_avalon_anti_slave_0_readdata;                                       // audio:fifo_full_s1_readdata -> audio_fifo_full_s1_translator:av_readdata
	wire    [1:0] audio_fifo_used_s1_translator_avalon_anti_slave_0_address;                                        // audio_fifo_used_s1_translator:av_address -> audio:fifo_used_s1_address
	wire   [31:0] audio_fifo_used_s1_translator_avalon_anti_slave_0_readdata;                                       // audio:fifo_used_s1_readdata -> audio_fifo_used_s1_translator:av_readdata
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest;                                 // cpu:jtag_debug_module_waitrequest -> cpu_jtag_debug_module_translator:av_waitrequest
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                   // cpu_jtag_debug_module_translator:av_writedata -> cpu:jtag_debug_module_writedata
	wire    [8:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_address;                                     // cpu_jtag_debug_module_translator:av_address -> cpu:jtag_debug_module_address
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_write;                                       // cpu_jtag_debug_module_translator:av_write -> cpu:jtag_debug_module_write
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_read;                                        // cpu_jtag_debug_module_translator:av_read -> cpu:jtag_debug_module_read
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                    // cpu:jtag_debug_module_readdata -> cpu_jtag_debug_module_translator:av_readdata
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                 // cpu_jtag_debug_module_translator:av_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire    [3:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                  // cpu_jtag_debug_module_translator:av_byteenable -> cpu:jtag_debug_module_byteenable
	wire   [31:0] audio_out_data_audio_s1_translator_avalon_anti_slave_0_writedata;                                 // audio_out_data_audio_s1_translator:av_writedata -> audio:out_data_audio_s1_writedata
	wire    [1:0] audio_out_data_audio_s1_translator_avalon_anti_slave_0_address;                                   // audio_out_data_audio_s1_translator:av_address -> audio:out_data_audio_s1_address
	wire          audio_out_data_audio_s1_translator_avalon_anti_slave_0_chipselect;                                // audio_out_data_audio_s1_translator:av_chipselect -> audio:out_data_audio_s1_chipselect
	wire          audio_out_data_audio_s1_translator_avalon_anti_slave_0_write;                                     // audio_out_data_audio_s1_translator:av_write -> audio:out_data_audio_s1_write_n
	wire   [31:0] audio_out_data_audio_s1_translator_avalon_anti_slave_0_readdata;                                  // audio:out_data_audio_s1_readdata -> audio_out_data_audio_s1_translator:av_readdata
	wire   [31:0] audio_out_pause_s1_translator_avalon_anti_slave_0_writedata;                                      // audio_out_pause_s1_translator:av_writedata -> audio:out_pause_s1_writedata
	wire    [1:0] audio_out_pause_s1_translator_avalon_anti_slave_0_address;                                        // audio_out_pause_s1_translator:av_address -> audio:out_pause_s1_address
	wire          audio_out_pause_s1_translator_avalon_anti_slave_0_chipselect;                                     // audio_out_pause_s1_translator:av_chipselect -> audio:out_pause_s1_chipselect
	wire          audio_out_pause_s1_translator_avalon_anti_slave_0_write;                                          // audio_out_pause_s1_translator:av_write -> audio:out_pause_s1_write_n
	wire   [31:0] audio_out_pause_s1_translator_avalon_anti_slave_0_readdata;                                       // audio:out_pause_s1_readdata -> audio_out_pause_s1_translator:av_readdata
	wire   [31:0] audio_out_stop_s1_translator_avalon_anti_slave_0_writedata;                                       // audio_out_stop_s1_translator:av_writedata -> audio:out_stop_s1_writedata
	wire    [1:0] audio_out_stop_s1_translator_avalon_anti_slave_0_address;                                         // audio_out_stop_s1_translator:av_address -> audio:out_stop_s1_address
	wire          audio_out_stop_s1_translator_avalon_anti_slave_0_chipselect;                                      // audio_out_stop_s1_translator:av_chipselect -> audio:out_stop_s1_chipselect
	wire          audio_out_stop_s1_translator_avalon_anti_slave_0_write;                                           // audio_out_stop_s1_translator:av_write -> audio:out_stop_s1_write_n
	wire   [31:0] audio_out_stop_s1_translator_avalon_anti_slave_0_readdata;                                        // audio:out_stop_s1_readdata -> audio_out_stop_s1_translator:av_readdata
	wire   [15:0] timer_s1_translator_avalon_anti_slave_0_writedata;                                                // timer_s1_translator:av_writedata -> timer:writedata
	wire    [2:0] timer_s1_translator_avalon_anti_slave_0_address;                                                  // timer_s1_translator:av_address -> timer:address
	wire          timer_s1_translator_avalon_anti_slave_0_chipselect;                                               // timer_s1_translator:av_chipselect -> timer:chipselect
	wire          timer_s1_translator_avalon_anti_slave_0_write;                                                    // timer_s1_translator:av_write -> timer:write_n
	wire   [15:0] timer_s1_translator_avalon_anti_slave_0_readdata;                                                 // timer:readdata -> timer_s1_translator:av_readdata
	wire   [31:0] key_s1_translator_avalon_anti_slave_0_writedata;                                                  // key_s1_translator:av_writedata -> key:writedata
	wire    [1:0] key_s1_translator_avalon_anti_slave_0_address;                                                    // key_s1_translator:av_address -> key:address
	wire          key_s1_translator_avalon_anti_slave_0_chipselect;                                                 // key_s1_translator:av_chipselect -> key:chipselect
	wire          key_s1_translator_avalon_anti_slave_0_write;                                                      // key_s1_translator:av_write -> key:write_n
	wire   [31:0] key_s1_translator_avalon_anti_slave_0_readdata;                                                   // key:readdata -> key_s1_translator:av_readdata
	wire   [31:0] signal_selector_s1_translator_avalon_anti_slave_0_writedata;                                      // signal_selector_s1_translator:av_writedata -> signal_selector:writedata
	wire    [1:0] signal_selector_s1_translator_avalon_anti_slave_0_address;                                        // signal_selector_s1_translator:av_address -> signal_selector:address
	wire          signal_selector_s1_translator_avalon_anti_slave_0_chipselect;                                     // signal_selector_s1_translator:av_chipselect -> signal_selector:chipselect
	wire          signal_selector_s1_translator_avalon_anti_slave_0_write;                                          // signal_selector_s1_translator:av_write -> signal_selector:write_n
	wire   [31:0] signal_selector_s1_translator_avalon_anti_slave_0_readdata;                                       // signal_selector:readdata -> signal_selector_s1_translator:av_readdata
	wire   [31:0] modulation_selector_s1_translator_avalon_anti_slave_0_writedata;                                  // modulation_selector_s1_translator:av_writedata -> modulation_selector:writedata
	wire    [1:0] modulation_selector_s1_translator_avalon_anti_slave_0_address;                                    // modulation_selector_s1_translator:av_address -> modulation_selector:address
	wire          modulation_selector_s1_translator_avalon_anti_slave_0_chipselect;                                 // modulation_selector_s1_translator:av_chipselect -> modulation_selector:chipselect
	wire          modulation_selector_s1_translator_avalon_anti_slave_0_write;                                      // modulation_selector_s1_translator:av_write -> modulation_selector:write_n
	wire   [31:0] modulation_selector_s1_translator_avalon_anti_slave_0_readdata;                                   // modulation_selector:readdata -> modulation_selector_s1_translator:av_readdata
	wire    [1:0] keyboard_keys_s1_translator_avalon_anti_slave_0_address;                                          // keyboard_keys_s1_translator:av_address -> keyboard_keys:address
	wire   [31:0] keyboard_keys_s1_translator_avalon_anti_slave_0_readdata;                                         // keyboard_keys:readdata -> keyboard_keys_s1_translator:av_readdata
	wire    [1:0] mouse_pos_s1_translator_avalon_anti_slave_0_address;                                              // mouse_pos_s1_translator:av_address -> mouse_pos:address
	wire   [31:0] mouse_pos_s1_translator_avalon_anti_slave_0_readdata;                                             // mouse_pos:readdata -> mouse_pos_s1_translator:av_readdata
	wire   [31:0] div_freq_s1_translator_avalon_anti_slave_0_writedata;                                             // div_freq_s1_translator:av_writedata -> div_freq:writedata
	wire    [1:0] div_freq_s1_translator_avalon_anti_slave_0_address;                                               // div_freq_s1_translator:av_address -> div_freq:address
	wire          div_freq_s1_translator_avalon_anti_slave_0_chipselect;                                            // div_freq_s1_translator:av_chipselect -> div_freq:chipselect
	wire          div_freq_s1_translator_avalon_anti_slave_0_write;                                                 // div_freq_s1_translator:av_write -> div_freq:write_n
	wire   [31:0] div_freq_s1_translator_avalon_anti_slave_0_readdata;                                              // div_freq:readdata -> div_freq_s1_translator:av_readdata
	wire   [31:0] audio_sel_s1_translator_avalon_anti_slave_0_writedata;                                            // audio_sel_s1_translator:av_writedata -> audio_sel:writedata
	wire    [1:0] audio_sel_s1_translator_avalon_anti_slave_0_address;                                              // audio_sel_s1_translator:av_address -> audio_sel:address
	wire          audio_sel_s1_translator_avalon_anti_slave_0_chipselect;                                           // audio_sel_s1_translator:av_chipselect -> audio_sel:chipselect
	wire          audio_sel_s1_translator_avalon_anti_slave_0_write;                                                // audio_sel_s1_translator:av_write -> audio_sel:write_n
	wire   [31:0] audio_sel_s1_translator_avalon_anti_slave_0_readdata;                                             // audio_sel:readdata -> audio_sel_s1_translator:av_readdata
	wire   [31:0] vga_to_nios_2_datamaster_translator_avalon_anti_slave_0_writedata;                                // vga_to_nios_2_datamaster_translator:av_writedata -> vga:to_nios_2_datamaster_writedata
	wire    [4:0] vga_to_nios_2_datamaster_translator_avalon_anti_slave_0_address;                                  // vga_to_nios_2_datamaster_translator:av_address -> vga:to_nios_2_datamaster_address
	wire          vga_to_nios_2_datamaster_translator_avalon_anti_slave_0_write;                                    // vga_to_nios_2_datamaster_translator:av_write -> vga:to_nios_2_datamaster_write
	wire          vga_to_nios_2_datamaster_translator_avalon_anti_slave_0_read;                                     // vga_to_nios_2_datamaster_translator:av_read -> vga:to_nios_2_datamaster_read
	wire   [31:0] vga_to_nios_2_datamaster_translator_avalon_anti_slave_0_readdata;                                 // vga:to_nios_2_datamaster_readdata -> vga_to_nios_2_datamaster_translator:av_readdata
	wire   [31:0] audio_wrclk_s1_translator_avalon_anti_slave_0_writedata;                                          // audio_wrclk_s1_translator:av_writedata -> audio:wrclk_s1_writedata
	wire    [1:0] audio_wrclk_s1_translator_avalon_anti_slave_0_address;                                            // audio_wrclk_s1_translator:av_address -> audio:wrclk_s1_address
	wire          audio_wrclk_s1_translator_avalon_anti_slave_0_chipselect;                                         // audio_wrclk_s1_translator:av_chipselect -> audio:wrclk_s1_chipselect
	wire          audio_wrclk_s1_translator_avalon_anti_slave_0_write;                                              // audio_wrclk_s1_translator:av_write -> audio:wrclk_s1_write_n
	wire   [31:0] audio_wrclk_s1_translator_avalon_anti_slave_0_readdata;                                           // audio:wrclk_s1_readdata -> audio_wrclk_s1_translator:av_readdata
	wire   [31:0] audio_wrreq_s1_translator_avalon_anti_slave_0_writedata;                                          // audio_wrreq_s1_translator:av_writedata -> audio:wrreq_s1_writedata
	wire    [1:0] audio_wrreq_s1_translator_avalon_anti_slave_0_address;                                            // audio_wrreq_s1_translator:av_address -> audio:wrreq_s1_address
	wire          audio_wrreq_s1_translator_avalon_anti_slave_0_chipselect;                                         // audio_wrreq_s1_translator:av_chipselect -> audio:wrreq_s1_chipselect
	wire          audio_wrreq_s1_translator_avalon_anti_slave_0_write;                                              // audio_wrreq_s1_translator:av_write -> audio:wrreq_s1_write_n
	wire   [31:0] audio_wrreq_s1_translator_avalon_anti_slave_0_readdata;                                           // audio:wrreq_s1_readdata -> audio_wrreq_s1_translator:av_readdata
	wire          sdram_s1_translator_avalon_anti_slave_0_waitrequest;                                              // sdram:za_waitrequest -> sdram_s1_translator:av_waitrequest
	wire   [15:0] sdram_s1_translator_avalon_anti_slave_0_writedata;                                                // sdram_s1_translator:av_writedata -> sdram:az_data
	wire   [21:0] sdram_s1_translator_avalon_anti_slave_0_address;                                                  // sdram_s1_translator:av_address -> sdram:az_addr
	wire          sdram_s1_translator_avalon_anti_slave_0_chipselect;                                               // sdram_s1_translator:av_chipselect -> sdram:az_cs
	wire          sdram_s1_translator_avalon_anti_slave_0_write;                                                    // sdram_s1_translator:av_write -> sdram:az_wr_n
	wire          sdram_s1_translator_avalon_anti_slave_0_read;                                                     // sdram_s1_translator:av_read -> sdram:az_rd_n
	wire   [15:0] sdram_s1_translator_avalon_anti_slave_0_readdata;                                                 // sdram:za_data -> sdram_s1_translator:av_readdata
	wire          sdram_s1_translator_avalon_anti_slave_0_readdatavalid;                                            // sdram:za_valid -> sdram_s1_translator:av_readdatavalid
	wire    [1:0] sdram_s1_translator_avalon_anti_slave_0_byteenable;                                               // sdram_s1_translator:av_byteenable -> sdram:az_be_n
	wire   [31:0] lfsr_clk_interrupt_gen_s1_translator_avalon_anti_slave_0_writedata;                               // lfsr_clk_interrupt_gen_s1_translator:av_writedata -> lfsr_clk_interrupt_gen:writedata
	wire    [1:0] lfsr_clk_interrupt_gen_s1_translator_avalon_anti_slave_0_address;                                 // lfsr_clk_interrupt_gen_s1_translator:av_address -> lfsr_clk_interrupt_gen:address
	wire          lfsr_clk_interrupt_gen_s1_translator_avalon_anti_slave_0_chipselect;                              // lfsr_clk_interrupt_gen_s1_translator:av_chipselect -> lfsr_clk_interrupt_gen:chipselect
	wire          lfsr_clk_interrupt_gen_s1_translator_avalon_anti_slave_0_write;                                   // lfsr_clk_interrupt_gen_s1_translator:av_write -> lfsr_clk_interrupt_gen:write_n
	wire   [31:0] lfsr_clk_interrupt_gen_s1_translator_avalon_anti_slave_0_readdata;                                // lfsr_clk_interrupt_gen:readdata -> lfsr_clk_interrupt_gen_s1_translator:av_readdata
	wire    [1:0] lfsr_val_s1_translator_avalon_anti_slave_0_address;                                               // lfsr_val_s1_translator:av_address -> lfsr_val:address
	wire   [31:0] lfsr_val_s1_translator_avalon_anti_slave_0_readdata;                                              // lfsr_val:readdata -> lfsr_val_s1_translator:av_readdata
	wire   [31:0] dds_increment_s1_translator_avalon_anti_slave_0_writedata;                                        // dds_increment_s1_translator:av_writedata -> dds_increment:writedata
	wire    [1:0] dds_increment_s1_translator_avalon_anti_slave_0_address;                                          // dds_increment_s1_translator:av_address -> dds_increment:address
	wire          dds_increment_s1_translator_avalon_anti_slave_0_chipselect;                                       // dds_increment_s1_translator:av_chipselect -> dds_increment:chipselect
	wire          dds_increment_s1_translator_avalon_anti_slave_0_write;                                            // dds_increment_s1_translator:av_write -> dds_increment:write_n
	wire   [31:0] dds_increment_s1_translator_avalon_anti_slave_0_readdata;                                         // dds_increment:readdata -> dds_increment_s1_translator:av_readdata
	wire          cpu_data_master_translator_avalon_universal_master_0_waitrequest;                                 // cpu_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_data_master_translator:uav_waitrequest
	wire    [2:0] cpu_data_master_translator_avalon_universal_master_0_burstcount;                                  // cpu_data_master_translator:uav_burstcount -> cpu_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_data_master_translator_avalon_universal_master_0_writedata;                                   // cpu_data_master_translator:uav_writedata -> cpu_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] cpu_data_master_translator_avalon_universal_master_0_address;                                     // cpu_data_master_translator:uav_address -> cpu_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_data_master_translator_avalon_universal_master_0_lock;                                        // cpu_data_master_translator:uav_lock -> cpu_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_data_master_translator_avalon_universal_master_0_write;                                       // cpu_data_master_translator:uav_write -> cpu_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_data_master_translator_avalon_universal_master_0_read;                                        // cpu_data_master_translator:uav_read -> cpu_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_data_master_translator_avalon_universal_master_0_readdata;                                    // cpu_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_data_master_translator:uav_readdata
	wire          cpu_data_master_translator_avalon_universal_master_0_debugaccess;                                 // cpu_data_master_translator:uav_debugaccess -> cpu_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_data_master_translator_avalon_universal_master_0_byteenable;                                  // cpu_data_master_translator:uav_byteenable -> cpu_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_data_master_translator_avalon_universal_master_0_readdatavalid;                               // cpu_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_data_master_translator:uav_readdatavalid
	wire          vga_to_sdram_translator_avalon_universal_master_0_waitrequest;                                    // vga_to_sdram_translator_avalon_universal_master_0_agent:av_waitrequest -> vga_to_sdram_translator:uav_waitrequest
	wire    [7:0] vga_to_sdram_translator_avalon_universal_master_0_burstcount;                                     // vga_to_sdram_translator:uav_burstcount -> vga_to_sdram_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] vga_to_sdram_translator_avalon_universal_master_0_writedata;                                      // vga_to_sdram_translator:uav_writedata -> vga_to_sdram_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] vga_to_sdram_translator_avalon_universal_master_0_address;                                        // vga_to_sdram_translator:uav_address -> vga_to_sdram_translator_avalon_universal_master_0_agent:av_address
	wire          vga_to_sdram_translator_avalon_universal_master_0_lock;                                           // vga_to_sdram_translator:uav_lock -> vga_to_sdram_translator_avalon_universal_master_0_agent:av_lock
	wire          vga_to_sdram_translator_avalon_universal_master_0_write;                                          // vga_to_sdram_translator:uav_write -> vga_to_sdram_translator_avalon_universal_master_0_agent:av_write
	wire          vga_to_sdram_translator_avalon_universal_master_0_read;                                           // vga_to_sdram_translator:uav_read -> vga_to_sdram_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] vga_to_sdram_translator_avalon_universal_master_0_readdata;                                       // vga_to_sdram_translator_avalon_universal_master_0_agent:av_readdata -> vga_to_sdram_translator:uav_readdata
	wire          vga_to_sdram_translator_avalon_universal_master_0_debugaccess;                                    // vga_to_sdram_translator:uav_debugaccess -> vga_to_sdram_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] vga_to_sdram_translator_avalon_universal_master_0_byteenable;                                     // vga_to_sdram_translator:uav_byteenable -> vga_to_sdram_translator_avalon_universal_master_0_agent:av_byteenable
	wire          vga_to_sdram_translator_avalon_universal_master_0_readdatavalid;                                  // vga_to_sdram_translator_avalon_universal_master_0_agent:av_readdatavalid -> vga_to_sdram_translator:uav_readdatavalid
	wire          cpu_instruction_master_translator_avalon_universal_master_0_waitrequest;                          // cpu_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_instruction_master_translator:uav_waitrequest
	wire    [2:0] cpu_instruction_master_translator_avalon_universal_master_0_burstcount;                           // cpu_instruction_master_translator:uav_burstcount -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_instruction_master_translator_avalon_universal_master_0_writedata;                            // cpu_instruction_master_translator:uav_writedata -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] cpu_instruction_master_translator_avalon_universal_master_0_address;                              // cpu_instruction_master_translator:uav_address -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_instruction_master_translator_avalon_universal_master_0_lock;                                 // cpu_instruction_master_translator:uav_lock -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_instruction_master_translator_avalon_universal_master_0_write;                                // cpu_instruction_master_translator:uav_write -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_instruction_master_translator_avalon_universal_master_0_read;                                 // cpu_instruction_master_translator:uav_read -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_instruction_master_translator_avalon_universal_master_0_readdata;                             // cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_instruction_master_translator:uav_readdata
	wire          cpu_instruction_master_translator_avalon_universal_master_0_debugaccess;                          // cpu_instruction_master_translator:uav_debugaccess -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_instruction_master_translator_avalon_universal_master_0_byteenable;                           // cpu_instruction_master_translator:uav_byteenable -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid;                        // cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_instruction_master_translator:uav_readdatavalid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // jtag_uart_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_avalon_jtag_slave_translator:uav_writedata
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // jtag_uart_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // jtag_uart_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [114:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [114:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;        // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                // sysid_qsys_control_slave_translator:uav_waitrequest -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                 // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_qsys_control_slave_translator:uav_burstcount
	wire   [31:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                  // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_qsys_control_slave_translator:uav_writedata
	wire   [31:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                    // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_qsys_control_slave_translator:uav_address
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                      // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_qsys_control_slave_translator:uav_write
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                       // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_qsys_control_slave_translator:uav_lock
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                       // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_qsys_control_slave_translator:uav_read
	wire   [31:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                   // sysid_qsys_control_slave_translator:uav_readdata -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;              // sysid_qsys_control_slave_translator:uav_readdatavalid -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_qsys_control_slave_translator:uav_debugaccess
	wire    [3:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                 // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_qsys_control_slave_translator:uav_byteenable
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;         // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;               // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;       // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [114:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;               // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;      // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;            // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;    // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [114:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;             // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;            // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;          // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;           // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;          // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;          // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;           // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;          // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                    // audio_data_fregen_s1_translator:uav_waitrequest -> audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                     // audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> audio_data_fregen_s1_translator:uav_burstcount
	wire   [31:0] audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                      // audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> audio_data_fregen_s1_translator:uav_writedata
	wire   [31:0] audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_m0_address;                        // audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:m0_address -> audio_data_fregen_s1_translator:uav_address
	wire          audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_m0_write;                          // audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:m0_write -> audio_data_fregen_s1_translator:uav_write
	wire          audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_m0_lock;                           // audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:m0_lock -> audio_data_fregen_s1_translator:uav_lock
	wire          audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_m0_read;                           // audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:m0_read -> audio_data_fregen_s1_translator:uav_read
	wire   [31:0] audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                       // audio_data_fregen_s1_translator:uav_readdata -> audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                  // audio_data_fregen_s1_translator:uav_readdatavalid -> audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                    // audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> audio_data_fregen_s1_translator:uav_debugaccess
	wire    [3:0] audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                     // audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> audio_data_fregen_s1_translator:uav_byteenable
	wire          audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;             // audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                   // audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;           // audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [114:0] audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                    // audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                   // audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;          // audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                // audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;        // audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [114:0] audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                 // audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                // audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;              // audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;               // audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;              // audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;              // audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;               // audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;              // audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          audio_empty_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                          // audio_empty_s1_translator:uav_waitrequest -> audio_empty_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] audio_empty_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                           // audio_empty_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> audio_empty_s1_translator:uav_burstcount
	wire   [31:0] audio_empty_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                            // audio_empty_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> audio_empty_s1_translator:uav_writedata
	wire   [31:0] audio_empty_s1_translator_avalon_universal_slave_0_agent_m0_address;                              // audio_empty_s1_translator_avalon_universal_slave_0_agent:m0_address -> audio_empty_s1_translator:uav_address
	wire          audio_empty_s1_translator_avalon_universal_slave_0_agent_m0_write;                                // audio_empty_s1_translator_avalon_universal_slave_0_agent:m0_write -> audio_empty_s1_translator:uav_write
	wire          audio_empty_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                 // audio_empty_s1_translator_avalon_universal_slave_0_agent:m0_lock -> audio_empty_s1_translator:uav_lock
	wire          audio_empty_s1_translator_avalon_universal_slave_0_agent_m0_read;                                 // audio_empty_s1_translator_avalon_universal_slave_0_agent:m0_read -> audio_empty_s1_translator:uav_read
	wire   [31:0] audio_empty_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                             // audio_empty_s1_translator:uav_readdata -> audio_empty_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          audio_empty_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                        // audio_empty_s1_translator:uav_readdatavalid -> audio_empty_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          audio_empty_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                          // audio_empty_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> audio_empty_s1_translator:uav_debugaccess
	wire    [3:0] audio_empty_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                           // audio_empty_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> audio_empty_s1_translator:uav_byteenable
	wire          audio_empty_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                   // audio_empty_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> audio_empty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          audio_empty_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                         // audio_empty_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> audio_empty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          audio_empty_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                 // audio_empty_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> audio_empty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [114:0] audio_empty_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                          // audio_empty_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> audio_empty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          audio_empty_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                         // audio_empty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> audio_empty_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          audio_empty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                // audio_empty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> audio_empty_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          audio_empty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                      // audio_empty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> audio_empty_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          audio_empty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;              // audio_empty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> audio_empty_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [114:0] audio_empty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                       // audio_empty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> audio_empty_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          audio_empty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                      // audio_empty_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> audio_empty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          audio_empty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                    // audio_empty_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> audio_empty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] audio_empty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                     // audio_empty_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> audio_empty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          audio_empty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                    // audio_empty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> audio_empty_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          audio_empty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                    // audio_empty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> audio_empty_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] audio_empty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                     // audio_empty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> audio_empty_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          audio_empty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                    // audio_empty_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> audio_empty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // audio_fifo_full_s1_translator:uav_waitrequest -> audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> audio_fifo_full_s1_translator:uav_burstcount
	wire   [31:0] audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                        // audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> audio_fifo_full_s1_translator:uav_writedata
	wire   [31:0] audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_m0_address;                          // audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:m0_address -> audio_fifo_full_s1_translator:uav_address
	wire          audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_m0_write;                            // audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:m0_write -> audio_fifo_full_s1_translator:uav_write
	wire          audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_m0_lock;                             // audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:m0_lock -> audio_fifo_full_s1_translator:uav_lock
	wire          audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_m0_read;                             // audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:m0_read -> audio_fifo_full_s1_translator:uav_read
	wire   [31:0] audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                         // audio_fifo_full_s1_translator:uav_readdata -> audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // audio_fifo_full_s1_translator:uav_readdatavalid -> audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> audio_fifo_full_s1_translator:uav_debugaccess
	wire    [3:0] audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> audio_fifo_full_s1_translator:uav_byteenable
	wire          audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [114:0] audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                      // audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [114:0] audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                // audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                 // audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                // audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // audio_fifo_used_s1_translator:uav_waitrequest -> audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> audio_fifo_used_s1_translator:uav_burstcount
	wire   [31:0] audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                        // audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> audio_fifo_used_s1_translator:uav_writedata
	wire   [31:0] audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_m0_address;                          // audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:m0_address -> audio_fifo_used_s1_translator:uav_address
	wire          audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_m0_write;                            // audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:m0_write -> audio_fifo_used_s1_translator:uav_write
	wire          audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_m0_lock;                             // audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:m0_lock -> audio_fifo_used_s1_translator:uav_lock
	wire          audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_m0_read;                             // audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:m0_read -> audio_fifo_used_s1_translator:uav_read
	wire   [31:0] audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                         // audio_fifo_used_s1_translator:uav_readdata -> audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // audio_fifo_used_s1_translator:uav_readdatavalid -> audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> audio_fifo_used_s1_translator:uav_debugaccess
	wire    [3:0] audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> audio_fifo_used_s1_translator:uav_byteenable
	wire          audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [114:0] audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                      // audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [114:0] audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                // audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                 // audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                // audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // cpu_jtag_debug_module_translator:uav_waitrequest -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                     // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_jtag_debug_module_translator:uav_writedata
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                       // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu_jtag_debug_module_translator:uav_address
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                         // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu_jtag_debug_module_translator:uav_write
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                          // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_jtag_debug_module_translator:uav_lock
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                          // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu_jtag_debug_module_translator:uav_read
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                      // cpu_jtag_debug_module_translator:uav_readdata -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // cpu_jtag_debug_module_translator:uav_readdatavalid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_jtag_debug_module_translator:uav_byteenable
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [114:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                   // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [114:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;             // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;              // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;             // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                 // audio_out_data_audio_s1_translator:uav_waitrequest -> audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                  // audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> audio_out_data_audio_s1_translator:uav_burstcount
	wire   [31:0] audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                   // audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> audio_out_data_audio_s1_translator:uav_writedata
	wire   [31:0] audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_m0_address;                     // audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:m0_address -> audio_out_data_audio_s1_translator:uav_address
	wire          audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_m0_write;                       // audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:m0_write -> audio_out_data_audio_s1_translator:uav_write
	wire          audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_m0_lock;                        // audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:m0_lock -> audio_out_data_audio_s1_translator:uav_lock
	wire          audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_m0_read;                        // audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:m0_read -> audio_out_data_audio_s1_translator:uav_read
	wire   [31:0] audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                    // audio_out_data_audio_s1_translator:uav_readdata -> audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;               // audio_out_data_audio_s1_translator:uav_readdatavalid -> audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                 // audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> audio_out_data_audio_s1_translator:uav_debugaccess
	wire    [3:0] audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                  // audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> audio_out_data_audio_s1_translator:uav_byteenable
	wire          audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;          // audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                // audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;        // audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [114:0] audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                 // audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                // audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;       // audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;             // audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;     // audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [114:0] audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;              // audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;             // audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;           // audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;            // audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;           // audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;           // audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;            // audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;           // audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          audio_out_pause_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // audio_out_pause_s1_translator:uav_waitrequest -> audio_out_pause_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] audio_out_pause_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // audio_out_pause_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> audio_out_pause_s1_translator:uav_burstcount
	wire   [31:0] audio_out_pause_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                        // audio_out_pause_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> audio_out_pause_s1_translator:uav_writedata
	wire   [31:0] audio_out_pause_s1_translator_avalon_universal_slave_0_agent_m0_address;                          // audio_out_pause_s1_translator_avalon_universal_slave_0_agent:m0_address -> audio_out_pause_s1_translator:uav_address
	wire          audio_out_pause_s1_translator_avalon_universal_slave_0_agent_m0_write;                            // audio_out_pause_s1_translator_avalon_universal_slave_0_agent:m0_write -> audio_out_pause_s1_translator:uav_write
	wire          audio_out_pause_s1_translator_avalon_universal_slave_0_agent_m0_lock;                             // audio_out_pause_s1_translator_avalon_universal_slave_0_agent:m0_lock -> audio_out_pause_s1_translator:uav_lock
	wire          audio_out_pause_s1_translator_avalon_universal_slave_0_agent_m0_read;                             // audio_out_pause_s1_translator_avalon_universal_slave_0_agent:m0_read -> audio_out_pause_s1_translator:uav_read
	wire   [31:0] audio_out_pause_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                         // audio_out_pause_s1_translator:uav_readdata -> audio_out_pause_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          audio_out_pause_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // audio_out_pause_s1_translator:uav_readdatavalid -> audio_out_pause_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          audio_out_pause_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // audio_out_pause_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> audio_out_pause_s1_translator:uav_debugaccess
	wire    [3:0] audio_out_pause_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // audio_out_pause_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> audio_out_pause_s1_translator:uav_byteenable
	wire          audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // audio_out_pause_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // audio_out_pause_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // audio_out_pause_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [114:0] audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                      // audio_out_pause_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> audio_out_pause_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> audio_out_pause_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> audio_out_pause_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> audio_out_pause_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [114:0] audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> audio_out_pause_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // audio_out_pause_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // audio_out_pause_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // audio_out_pause_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> audio_out_pause_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                // audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> audio_out_pause_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                 // audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> audio_out_pause_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                // audio_out_pause_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          audio_out_stop_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // audio_out_stop_s1_translator:uav_waitrequest -> audio_out_stop_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] audio_out_stop_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // audio_out_stop_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> audio_out_stop_s1_translator:uav_burstcount
	wire   [31:0] audio_out_stop_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                         // audio_out_stop_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> audio_out_stop_s1_translator:uav_writedata
	wire   [31:0] audio_out_stop_s1_translator_avalon_universal_slave_0_agent_m0_address;                           // audio_out_stop_s1_translator_avalon_universal_slave_0_agent:m0_address -> audio_out_stop_s1_translator:uav_address
	wire          audio_out_stop_s1_translator_avalon_universal_slave_0_agent_m0_write;                             // audio_out_stop_s1_translator_avalon_universal_slave_0_agent:m0_write -> audio_out_stop_s1_translator:uav_write
	wire          audio_out_stop_s1_translator_avalon_universal_slave_0_agent_m0_lock;                              // audio_out_stop_s1_translator_avalon_universal_slave_0_agent:m0_lock -> audio_out_stop_s1_translator:uav_lock
	wire          audio_out_stop_s1_translator_avalon_universal_slave_0_agent_m0_read;                              // audio_out_stop_s1_translator_avalon_universal_slave_0_agent:m0_read -> audio_out_stop_s1_translator:uav_read
	wire   [31:0] audio_out_stop_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                          // audio_out_stop_s1_translator:uav_readdata -> audio_out_stop_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          audio_out_stop_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // audio_out_stop_s1_translator:uav_readdatavalid -> audio_out_stop_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          audio_out_stop_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // audio_out_stop_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> audio_out_stop_s1_translator:uav_debugaccess
	wire    [3:0] audio_out_stop_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // audio_out_stop_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> audio_out_stop_s1_translator:uav_byteenable
	wire          audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // audio_out_stop_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // audio_out_stop_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // audio_out_stop_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [114:0] audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                       // audio_out_stop_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> audio_out_stop_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> audio_out_stop_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> audio_out_stop_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> audio_out_stop_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [114:0] audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> audio_out_stop_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // audio_out_stop_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // audio_out_stop_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // audio_out_stop_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> audio_out_stop_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                 // audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> audio_out_stop_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                  // audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> audio_out_stop_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                 // audio_out_stop_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // timer_s1_translator:uav_waitrequest -> timer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // timer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_s1_translator:uav_burstcount
	wire   [31:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // timer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_s1_translator:uav_writedata
	wire   [31:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // timer_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_s1_translator:uav_address
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // timer_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_s1_translator:uav_write
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // timer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_s1_translator:uav_lock
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // timer_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_s1_translator:uav_read
	wire   [31:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // timer_s1_translator:uav_readdata -> timer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // timer_s1_translator:uav_readdatavalid -> timer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // timer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_s1_translator:uav_debugaccess
	wire    [3:0] timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // timer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_s1_translator:uav_byteenable
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [114:0] timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // timer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [114:0] timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                          // timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                           // timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                          // timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          key_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // key_s1_translator:uav_waitrequest -> key_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] key_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // key_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> key_s1_translator:uav_burstcount
	wire   [31:0] key_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // key_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> key_s1_translator:uav_writedata
	wire   [31:0] key_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // key_s1_translator_avalon_universal_slave_0_agent:m0_address -> key_s1_translator:uav_address
	wire          key_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // key_s1_translator_avalon_universal_slave_0_agent:m0_write -> key_s1_translator:uav_write
	wire          key_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // key_s1_translator_avalon_universal_slave_0_agent:m0_lock -> key_s1_translator:uav_lock
	wire          key_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // key_s1_translator_avalon_universal_slave_0_agent:m0_read -> key_s1_translator:uav_read
	wire   [31:0] key_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // key_s1_translator:uav_readdata -> key_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          key_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // key_s1_translator:uav_readdatavalid -> key_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          key_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // key_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> key_s1_translator:uav_debugaccess
	wire    [3:0] key_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // key_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> key_s1_translator:uav_byteenable
	wire          key_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // key_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          key_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // key_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          key_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // key_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [114:0] key_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // key_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          key_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> key_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> key_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> key_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> key_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [114:0] key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> key_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // key_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                            // key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                             // key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                            // key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          signal_selector_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // signal_selector_s1_translator:uav_waitrequest -> signal_selector_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] signal_selector_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // signal_selector_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> signal_selector_s1_translator:uav_burstcount
	wire   [31:0] signal_selector_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                        // signal_selector_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> signal_selector_s1_translator:uav_writedata
	wire   [31:0] signal_selector_s1_translator_avalon_universal_slave_0_agent_m0_address;                          // signal_selector_s1_translator_avalon_universal_slave_0_agent:m0_address -> signal_selector_s1_translator:uav_address
	wire          signal_selector_s1_translator_avalon_universal_slave_0_agent_m0_write;                            // signal_selector_s1_translator_avalon_universal_slave_0_agent:m0_write -> signal_selector_s1_translator:uav_write
	wire          signal_selector_s1_translator_avalon_universal_slave_0_agent_m0_lock;                             // signal_selector_s1_translator_avalon_universal_slave_0_agent:m0_lock -> signal_selector_s1_translator:uav_lock
	wire          signal_selector_s1_translator_avalon_universal_slave_0_agent_m0_read;                             // signal_selector_s1_translator_avalon_universal_slave_0_agent:m0_read -> signal_selector_s1_translator:uav_read
	wire   [31:0] signal_selector_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                         // signal_selector_s1_translator:uav_readdata -> signal_selector_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          signal_selector_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // signal_selector_s1_translator:uav_readdatavalid -> signal_selector_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          signal_selector_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // signal_selector_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> signal_selector_s1_translator:uav_debugaccess
	wire    [3:0] signal_selector_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // signal_selector_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> signal_selector_s1_translator:uav_byteenable
	wire          signal_selector_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // signal_selector_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> signal_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          signal_selector_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // signal_selector_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> signal_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          signal_selector_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // signal_selector_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> signal_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [114:0] signal_selector_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                      // signal_selector_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> signal_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          signal_selector_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // signal_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> signal_selector_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          signal_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // signal_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> signal_selector_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          signal_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // signal_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> signal_selector_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          signal_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // signal_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> signal_selector_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [114:0] signal_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // signal_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> signal_selector_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          signal_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // signal_selector_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> signal_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          signal_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // signal_selector_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> signal_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] signal_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // signal_selector_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> signal_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          signal_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // signal_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> signal_selector_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          signal_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                // signal_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> signal_selector_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] signal_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                 // signal_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> signal_selector_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          signal_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                // signal_selector_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> signal_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          modulation_selector_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                  // modulation_selector_s1_translator:uav_waitrequest -> modulation_selector_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] modulation_selector_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                   // modulation_selector_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> modulation_selector_s1_translator:uav_burstcount
	wire   [31:0] modulation_selector_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                    // modulation_selector_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> modulation_selector_s1_translator:uav_writedata
	wire   [31:0] modulation_selector_s1_translator_avalon_universal_slave_0_agent_m0_address;                      // modulation_selector_s1_translator_avalon_universal_slave_0_agent:m0_address -> modulation_selector_s1_translator:uav_address
	wire          modulation_selector_s1_translator_avalon_universal_slave_0_agent_m0_write;                        // modulation_selector_s1_translator_avalon_universal_slave_0_agent:m0_write -> modulation_selector_s1_translator:uav_write
	wire          modulation_selector_s1_translator_avalon_universal_slave_0_agent_m0_lock;                         // modulation_selector_s1_translator_avalon_universal_slave_0_agent:m0_lock -> modulation_selector_s1_translator:uav_lock
	wire          modulation_selector_s1_translator_avalon_universal_slave_0_agent_m0_read;                         // modulation_selector_s1_translator_avalon_universal_slave_0_agent:m0_read -> modulation_selector_s1_translator:uav_read
	wire   [31:0] modulation_selector_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                     // modulation_selector_s1_translator:uav_readdata -> modulation_selector_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          modulation_selector_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                // modulation_selector_s1_translator:uav_readdatavalid -> modulation_selector_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          modulation_selector_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                  // modulation_selector_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> modulation_selector_s1_translator:uav_debugaccess
	wire    [3:0] modulation_selector_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                   // modulation_selector_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> modulation_selector_s1_translator:uav_byteenable
	wire          modulation_selector_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;           // modulation_selector_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> modulation_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          modulation_selector_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                 // modulation_selector_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> modulation_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          modulation_selector_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;         // modulation_selector_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> modulation_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [114:0] modulation_selector_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                  // modulation_selector_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> modulation_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          modulation_selector_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                 // modulation_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> modulation_selector_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          modulation_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;        // modulation_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> modulation_selector_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          modulation_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;              // modulation_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> modulation_selector_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          modulation_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;      // modulation_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> modulation_selector_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [114:0] modulation_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;               // modulation_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> modulation_selector_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          modulation_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;              // modulation_selector_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> modulation_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          modulation_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;            // modulation_selector_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> modulation_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] modulation_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;             // modulation_selector_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> modulation_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          modulation_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;            // modulation_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> modulation_selector_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          modulation_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;            // modulation_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> modulation_selector_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] modulation_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;             // modulation_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> modulation_selector_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          modulation_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;            // modulation_selector_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> modulation_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          keyboard_keys_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // keyboard_keys_s1_translator:uav_waitrequest -> keyboard_keys_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] keyboard_keys_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // keyboard_keys_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> keyboard_keys_s1_translator:uav_burstcount
	wire   [31:0] keyboard_keys_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                          // keyboard_keys_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> keyboard_keys_s1_translator:uav_writedata
	wire   [31:0] keyboard_keys_s1_translator_avalon_universal_slave_0_agent_m0_address;                            // keyboard_keys_s1_translator_avalon_universal_slave_0_agent:m0_address -> keyboard_keys_s1_translator:uav_address
	wire          keyboard_keys_s1_translator_avalon_universal_slave_0_agent_m0_write;                              // keyboard_keys_s1_translator_avalon_universal_slave_0_agent:m0_write -> keyboard_keys_s1_translator:uav_write
	wire          keyboard_keys_s1_translator_avalon_universal_slave_0_agent_m0_lock;                               // keyboard_keys_s1_translator_avalon_universal_slave_0_agent:m0_lock -> keyboard_keys_s1_translator:uav_lock
	wire          keyboard_keys_s1_translator_avalon_universal_slave_0_agent_m0_read;                               // keyboard_keys_s1_translator_avalon_universal_slave_0_agent:m0_read -> keyboard_keys_s1_translator:uav_read
	wire   [31:0] keyboard_keys_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                           // keyboard_keys_s1_translator:uav_readdata -> keyboard_keys_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          keyboard_keys_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // keyboard_keys_s1_translator:uav_readdatavalid -> keyboard_keys_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          keyboard_keys_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // keyboard_keys_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> keyboard_keys_s1_translator:uav_debugaccess
	wire    [3:0] keyboard_keys_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // keyboard_keys_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> keyboard_keys_s1_translator:uav_byteenable
	wire          keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // keyboard_keys_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // keyboard_keys_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // keyboard_keys_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [114:0] keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                        // keyboard_keys_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> keyboard_keys_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> keyboard_keys_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> keyboard_keys_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> keyboard_keys_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [114:0] keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> keyboard_keys_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // keyboard_keys_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // keyboard_keys_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // keyboard_keys_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> keyboard_keys_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                  // keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> keyboard_keys_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                   // keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> keyboard_keys_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                  // keyboard_keys_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          mouse_pos_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // mouse_pos_s1_translator:uav_waitrequest -> mouse_pos_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] mouse_pos_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // mouse_pos_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> mouse_pos_s1_translator:uav_burstcount
	wire   [31:0] mouse_pos_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // mouse_pos_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> mouse_pos_s1_translator:uav_writedata
	wire   [31:0] mouse_pos_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // mouse_pos_s1_translator_avalon_universal_slave_0_agent:m0_address -> mouse_pos_s1_translator:uav_address
	wire          mouse_pos_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // mouse_pos_s1_translator_avalon_universal_slave_0_agent:m0_write -> mouse_pos_s1_translator:uav_write
	wire          mouse_pos_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // mouse_pos_s1_translator_avalon_universal_slave_0_agent:m0_lock -> mouse_pos_s1_translator:uav_lock
	wire          mouse_pos_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // mouse_pos_s1_translator_avalon_universal_slave_0_agent:m0_read -> mouse_pos_s1_translator:uav_read
	wire   [31:0] mouse_pos_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // mouse_pos_s1_translator:uav_readdata -> mouse_pos_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          mouse_pos_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // mouse_pos_s1_translator:uav_readdatavalid -> mouse_pos_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          mouse_pos_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // mouse_pos_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> mouse_pos_s1_translator:uav_debugaccess
	wire    [3:0] mouse_pos_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // mouse_pos_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> mouse_pos_s1_translator:uav_byteenable
	wire          mouse_pos_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // mouse_pos_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> mouse_pos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          mouse_pos_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // mouse_pos_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> mouse_pos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          mouse_pos_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // mouse_pos_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> mouse_pos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [114:0] mouse_pos_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // mouse_pos_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> mouse_pos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          mouse_pos_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // mouse_pos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> mouse_pos_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          mouse_pos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // mouse_pos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> mouse_pos_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          mouse_pos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // mouse_pos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> mouse_pos_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          mouse_pos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // mouse_pos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> mouse_pos_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [114:0] mouse_pos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // mouse_pos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> mouse_pos_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          mouse_pos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // mouse_pos_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> mouse_pos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          mouse_pos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // mouse_pos_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> mouse_pos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] mouse_pos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // mouse_pos_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> mouse_pos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          mouse_pos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // mouse_pos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> mouse_pos_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          mouse_pos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                      // mouse_pos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> mouse_pos_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] mouse_pos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                       // mouse_pos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> mouse_pos_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          mouse_pos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                      // mouse_pos_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> mouse_pos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          div_freq_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // div_freq_s1_translator:uav_waitrequest -> div_freq_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] div_freq_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // div_freq_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> div_freq_s1_translator:uav_burstcount
	wire   [31:0] div_freq_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                               // div_freq_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> div_freq_s1_translator:uav_writedata
	wire   [31:0] div_freq_s1_translator_avalon_universal_slave_0_agent_m0_address;                                 // div_freq_s1_translator_avalon_universal_slave_0_agent:m0_address -> div_freq_s1_translator:uav_address
	wire          div_freq_s1_translator_avalon_universal_slave_0_agent_m0_write;                                   // div_freq_s1_translator_avalon_universal_slave_0_agent:m0_write -> div_freq_s1_translator:uav_write
	wire          div_freq_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                    // div_freq_s1_translator_avalon_universal_slave_0_agent:m0_lock -> div_freq_s1_translator:uav_lock
	wire          div_freq_s1_translator_avalon_universal_slave_0_agent_m0_read;                                    // div_freq_s1_translator_avalon_universal_slave_0_agent:m0_read -> div_freq_s1_translator:uav_read
	wire   [31:0] div_freq_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                // div_freq_s1_translator:uav_readdata -> div_freq_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          div_freq_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // div_freq_s1_translator:uav_readdatavalid -> div_freq_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          div_freq_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // div_freq_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> div_freq_s1_translator:uav_debugaccess
	wire    [3:0] div_freq_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // div_freq_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> div_freq_s1_translator:uav_byteenable
	wire          div_freq_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // div_freq_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> div_freq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          div_freq_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // div_freq_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> div_freq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          div_freq_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // div_freq_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> div_freq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [114:0] div_freq_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                             // div_freq_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> div_freq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          div_freq_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // div_freq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> div_freq_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          div_freq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // div_freq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> div_freq_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          div_freq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // div_freq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> div_freq_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          div_freq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // div_freq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> div_freq_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [114:0] div_freq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // div_freq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> div_freq_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          div_freq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // div_freq_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> div_freq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          div_freq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // div_freq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> div_freq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] div_freq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // div_freq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> div_freq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          div_freq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // div_freq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> div_freq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          div_freq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                       // div_freq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> div_freq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] div_freq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                        // div_freq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> div_freq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          div_freq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                       // div_freq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> div_freq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          audio_sel_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // audio_sel_s1_translator:uav_waitrequest -> audio_sel_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] audio_sel_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // audio_sel_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> audio_sel_s1_translator:uav_burstcount
	wire   [31:0] audio_sel_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // audio_sel_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> audio_sel_s1_translator:uav_writedata
	wire   [31:0] audio_sel_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // audio_sel_s1_translator_avalon_universal_slave_0_agent:m0_address -> audio_sel_s1_translator:uav_address
	wire          audio_sel_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // audio_sel_s1_translator_avalon_universal_slave_0_agent:m0_write -> audio_sel_s1_translator:uav_write
	wire          audio_sel_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // audio_sel_s1_translator_avalon_universal_slave_0_agent:m0_lock -> audio_sel_s1_translator:uav_lock
	wire          audio_sel_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // audio_sel_s1_translator_avalon_universal_slave_0_agent:m0_read -> audio_sel_s1_translator:uav_read
	wire   [31:0] audio_sel_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // audio_sel_s1_translator:uav_readdata -> audio_sel_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          audio_sel_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // audio_sel_s1_translator:uav_readdatavalid -> audio_sel_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          audio_sel_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // audio_sel_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> audio_sel_s1_translator:uav_debugaccess
	wire    [3:0] audio_sel_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // audio_sel_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> audio_sel_s1_translator:uav_byteenable
	wire          audio_sel_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // audio_sel_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> audio_sel_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          audio_sel_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // audio_sel_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> audio_sel_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          audio_sel_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // audio_sel_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> audio_sel_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [114:0] audio_sel_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // audio_sel_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> audio_sel_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          audio_sel_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // audio_sel_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> audio_sel_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          audio_sel_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // audio_sel_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> audio_sel_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          audio_sel_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // audio_sel_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> audio_sel_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          audio_sel_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // audio_sel_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> audio_sel_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [114:0] audio_sel_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // audio_sel_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> audio_sel_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          audio_sel_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // audio_sel_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> audio_sel_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          audio_sel_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // audio_sel_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> audio_sel_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] audio_sel_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // audio_sel_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> audio_sel_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          audio_sel_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // audio_sel_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> audio_sel_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          audio_sel_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                      // audio_sel_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> audio_sel_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] audio_sel_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                       // audio_sel_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> audio_sel_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          audio_sel_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                      // audio_sel_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> audio_sel_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_m0_waitrequest;                // vga_to_nios_2_datamaster_translator:uav_waitrequest -> vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_m0_burstcount;                 // vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:m0_burstcount -> vga_to_nios_2_datamaster_translator:uav_burstcount
	wire   [31:0] vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_m0_writedata;                  // vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:m0_writedata -> vga_to_nios_2_datamaster_translator:uav_writedata
	wire   [31:0] vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_m0_address;                    // vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:m0_address -> vga_to_nios_2_datamaster_translator:uav_address
	wire          vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_m0_write;                      // vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:m0_write -> vga_to_nios_2_datamaster_translator:uav_write
	wire          vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_m0_lock;                       // vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:m0_lock -> vga_to_nios_2_datamaster_translator:uav_lock
	wire          vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_m0_read;                       // vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:m0_read -> vga_to_nios_2_datamaster_translator:uav_read
	wire   [31:0] vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_m0_readdata;                   // vga_to_nios_2_datamaster_translator:uav_readdata -> vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_m0_readdatavalid;              // vga_to_nios_2_datamaster_translator:uav_readdatavalid -> vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_m0_debugaccess;                // vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:m0_debugaccess -> vga_to_nios_2_datamaster_translator:uav_debugaccess
	wire    [3:0] vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_m0_byteenable;                 // vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:m0_byteenable -> vga_to_nios_2_datamaster_translator:uav_byteenable
	wire          vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;         // vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rf_source_valid;               // vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:rf_source_valid -> vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;       // vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [114:0] vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rf_source_data;                // vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:rf_source_data -> vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rf_source_ready;               // vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;      // vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;            // vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;    // vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [114:0] vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;             // vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;            // vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:rf_sink_ready -> vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;          // vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;           // vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;          // vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;          // vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;           // vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;          // vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          audio_wrclk_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                          // audio_wrclk_s1_translator:uav_waitrequest -> audio_wrclk_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] audio_wrclk_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                           // audio_wrclk_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> audio_wrclk_s1_translator:uav_burstcount
	wire   [31:0] audio_wrclk_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                            // audio_wrclk_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> audio_wrclk_s1_translator:uav_writedata
	wire   [31:0] audio_wrclk_s1_translator_avalon_universal_slave_0_agent_m0_address;                              // audio_wrclk_s1_translator_avalon_universal_slave_0_agent:m0_address -> audio_wrclk_s1_translator:uav_address
	wire          audio_wrclk_s1_translator_avalon_universal_slave_0_agent_m0_write;                                // audio_wrclk_s1_translator_avalon_universal_slave_0_agent:m0_write -> audio_wrclk_s1_translator:uav_write
	wire          audio_wrclk_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                 // audio_wrclk_s1_translator_avalon_universal_slave_0_agent:m0_lock -> audio_wrclk_s1_translator:uav_lock
	wire          audio_wrclk_s1_translator_avalon_universal_slave_0_agent_m0_read;                                 // audio_wrclk_s1_translator_avalon_universal_slave_0_agent:m0_read -> audio_wrclk_s1_translator:uav_read
	wire   [31:0] audio_wrclk_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                             // audio_wrclk_s1_translator:uav_readdata -> audio_wrclk_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          audio_wrclk_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                        // audio_wrclk_s1_translator:uav_readdatavalid -> audio_wrclk_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          audio_wrclk_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                          // audio_wrclk_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> audio_wrclk_s1_translator:uav_debugaccess
	wire    [3:0] audio_wrclk_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                           // audio_wrclk_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> audio_wrclk_s1_translator:uav_byteenable
	wire          audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                   // audio_wrclk_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                         // audio_wrclk_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                 // audio_wrclk_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [114:0] audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                          // audio_wrclk_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                         // audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> audio_wrclk_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                // audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> audio_wrclk_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                      // audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> audio_wrclk_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;              // audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> audio_wrclk_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [114:0] audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                       // audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> audio_wrclk_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                      // audio_wrclk_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                    // audio_wrclk_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                     // audio_wrclk_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                    // audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> audio_wrclk_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                    // audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> audio_wrclk_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                     // audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> audio_wrclk_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                    // audio_wrclk_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          audio_wrreq_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                          // audio_wrreq_s1_translator:uav_waitrequest -> audio_wrreq_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] audio_wrreq_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                           // audio_wrreq_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> audio_wrreq_s1_translator:uav_burstcount
	wire   [31:0] audio_wrreq_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                            // audio_wrreq_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> audio_wrreq_s1_translator:uav_writedata
	wire   [31:0] audio_wrreq_s1_translator_avalon_universal_slave_0_agent_m0_address;                              // audio_wrreq_s1_translator_avalon_universal_slave_0_agent:m0_address -> audio_wrreq_s1_translator:uav_address
	wire          audio_wrreq_s1_translator_avalon_universal_slave_0_agent_m0_write;                                // audio_wrreq_s1_translator_avalon_universal_slave_0_agent:m0_write -> audio_wrreq_s1_translator:uav_write
	wire          audio_wrreq_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                 // audio_wrreq_s1_translator_avalon_universal_slave_0_agent:m0_lock -> audio_wrreq_s1_translator:uav_lock
	wire          audio_wrreq_s1_translator_avalon_universal_slave_0_agent_m0_read;                                 // audio_wrreq_s1_translator_avalon_universal_slave_0_agent:m0_read -> audio_wrreq_s1_translator:uav_read
	wire   [31:0] audio_wrreq_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                             // audio_wrreq_s1_translator:uav_readdata -> audio_wrreq_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          audio_wrreq_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                        // audio_wrreq_s1_translator:uav_readdatavalid -> audio_wrreq_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          audio_wrreq_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                          // audio_wrreq_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> audio_wrreq_s1_translator:uav_debugaccess
	wire    [3:0] audio_wrreq_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                           // audio_wrreq_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> audio_wrreq_s1_translator:uav_byteenable
	wire          audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                   // audio_wrreq_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                         // audio_wrreq_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                 // audio_wrreq_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [114:0] audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                          // audio_wrreq_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                         // audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> audio_wrreq_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                // audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> audio_wrreq_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                      // audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> audio_wrreq_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;              // audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> audio_wrreq_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [114:0] audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                       // audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> audio_wrreq_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                      // audio_wrreq_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                    // audio_wrreq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                     // audio_wrreq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                    // audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> audio_wrreq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                    // audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> audio_wrreq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                     // audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> audio_wrreq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                    // audio_wrreq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // sdram_s1_translator:uav_waitrequest -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // sdram_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_s1_translator:uav_burstcount
	wire   [15:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // sdram_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_s1_translator:uav_writedata
	wire   [31:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // sdram_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdram_s1_translator:uav_address
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // sdram_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdram_s1_translator:uav_write
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // sdram_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_s1_translator:uav_lock
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // sdram_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdram_s1_translator:uav_read
	wire   [15:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // sdram_s1_translator:uav_readdata -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // sdram_s1_translator:uav_readdatavalid -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // sdram_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_s1_translator:uav_debugaccess
	wire    [1:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // sdram_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_s1_translator:uav_byteenable
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [96:0] sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [96:0] sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [17:0] sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                          // sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [17:0] sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                           // sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                          // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;               // lfsr_clk_interrupt_gen_s1_translator:uav_waitrequest -> lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                // lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> lfsr_clk_interrupt_gen_s1_translator:uav_burstcount
	wire   [31:0] lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                 // lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> lfsr_clk_interrupt_gen_s1_translator:uav_writedata
	wire   [31:0] lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_m0_address;                   // lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:m0_address -> lfsr_clk_interrupt_gen_s1_translator:uav_address
	wire          lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_m0_write;                     // lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:m0_write -> lfsr_clk_interrupt_gen_s1_translator:uav_write
	wire          lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_m0_lock;                      // lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:m0_lock -> lfsr_clk_interrupt_gen_s1_translator:uav_lock
	wire          lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_m0_read;                      // lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:m0_read -> lfsr_clk_interrupt_gen_s1_translator:uav_read
	wire   [31:0] lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                  // lfsr_clk_interrupt_gen_s1_translator:uav_readdata -> lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;             // lfsr_clk_interrupt_gen_s1_translator:uav_readdatavalid -> lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;               // lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> lfsr_clk_interrupt_gen_s1_translator:uav_debugaccess
	wire    [3:0] lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                // lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> lfsr_clk_interrupt_gen_s1_translator:uav_byteenable
	wire          lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;        // lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;              // lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;      // lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [114:0] lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rf_source_data;               // lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;              // lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;     // lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;           // lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;   // lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [114:0] lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;            // lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;           // lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;         // lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;          // lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;         // lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;         // lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;          // lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;         // lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          lfsr_val_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // lfsr_val_s1_translator:uav_waitrequest -> lfsr_val_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] lfsr_val_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // lfsr_val_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> lfsr_val_s1_translator:uav_burstcount
	wire   [31:0] lfsr_val_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                               // lfsr_val_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> lfsr_val_s1_translator:uav_writedata
	wire   [31:0] lfsr_val_s1_translator_avalon_universal_slave_0_agent_m0_address;                                 // lfsr_val_s1_translator_avalon_universal_slave_0_agent:m0_address -> lfsr_val_s1_translator:uav_address
	wire          lfsr_val_s1_translator_avalon_universal_slave_0_agent_m0_write;                                   // lfsr_val_s1_translator_avalon_universal_slave_0_agent:m0_write -> lfsr_val_s1_translator:uav_write
	wire          lfsr_val_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                    // lfsr_val_s1_translator_avalon_universal_slave_0_agent:m0_lock -> lfsr_val_s1_translator:uav_lock
	wire          lfsr_val_s1_translator_avalon_universal_slave_0_agent_m0_read;                                    // lfsr_val_s1_translator_avalon_universal_slave_0_agent:m0_read -> lfsr_val_s1_translator:uav_read
	wire   [31:0] lfsr_val_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                // lfsr_val_s1_translator:uav_readdata -> lfsr_val_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          lfsr_val_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // lfsr_val_s1_translator:uav_readdatavalid -> lfsr_val_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          lfsr_val_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // lfsr_val_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> lfsr_val_s1_translator:uav_debugaccess
	wire    [3:0] lfsr_val_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // lfsr_val_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> lfsr_val_s1_translator:uav_byteenable
	wire          lfsr_val_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // lfsr_val_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> lfsr_val_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          lfsr_val_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // lfsr_val_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> lfsr_val_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          lfsr_val_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // lfsr_val_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> lfsr_val_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [114:0] lfsr_val_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                             // lfsr_val_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> lfsr_val_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          lfsr_val_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // lfsr_val_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> lfsr_val_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          lfsr_val_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // lfsr_val_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> lfsr_val_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          lfsr_val_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // lfsr_val_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> lfsr_val_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          lfsr_val_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // lfsr_val_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> lfsr_val_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [114:0] lfsr_val_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // lfsr_val_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> lfsr_val_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          lfsr_val_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // lfsr_val_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> lfsr_val_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          lfsr_val_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // lfsr_val_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> lfsr_val_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] lfsr_val_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // lfsr_val_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> lfsr_val_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          lfsr_val_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // lfsr_val_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> lfsr_val_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          lfsr_val_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                       // lfsr_val_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> lfsr_val_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] lfsr_val_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                        // lfsr_val_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> lfsr_val_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          lfsr_val_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                       // lfsr_val_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> lfsr_val_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          dds_increment_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // dds_increment_s1_translator:uav_waitrequest -> dds_increment_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] dds_increment_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // dds_increment_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> dds_increment_s1_translator:uav_burstcount
	wire   [31:0] dds_increment_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                          // dds_increment_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> dds_increment_s1_translator:uav_writedata
	wire   [31:0] dds_increment_s1_translator_avalon_universal_slave_0_agent_m0_address;                            // dds_increment_s1_translator_avalon_universal_slave_0_agent:m0_address -> dds_increment_s1_translator:uav_address
	wire          dds_increment_s1_translator_avalon_universal_slave_0_agent_m0_write;                              // dds_increment_s1_translator_avalon_universal_slave_0_agent:m0_write -> dds_increment_s1_translator:uav_write
	wire          dds_increment_s1_translator_avalon_universal_slave_0_agent_m0_lock;                               // dds_increment_s1_translator_avalon_universal_slave_0_agent:m0_lock -> dds_increment_s1_translator:uav_lock
	wire          dds_increment_s1_translator_avalon_universal_slave_0_agent_m0_read;                               // dds_increment_s1_translator_avalon_universal_slave_0_agent:m0_read -> dds_increment_s1_translator:uav_read
	wire   [31:0] dds_increment_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                           // dds_increment_s1_translator:uav_readdata -> dds_increment_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          dds_increment_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // dds_increment_s1_translator:uav_readdatavalid -> dds_increment_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          dds_increment_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // dds_increment_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> dds_increment_s1_translator:uav_debugaccess
	wire    [3:0] dds_increment_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // dds_increment_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> dds_increment_s1_translator:uav_byteenable
	wire          dds_increment_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // dds_increment_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> dds_increment_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          dds_increment_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // dds_increment_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> dds_increment_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          dds_increment_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // dds_increment_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> dds_increment_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [114:0] dds_increment_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                        // dds_increment_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> dds_increment_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          dds_increment_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // dds_increment_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> dds_increment_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          dds_increment_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // dds_increment_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> dds_increment_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          dds_increment_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // dds_increment_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> dds_increment_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          dds_increment_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // dds_increment_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> dds_increment_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [114:0] dds_increment_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // dds_increment_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> dds_increment_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          dds_increment_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // dds_increment_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> dds_increment_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          dds_increment_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // dds_increment_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> dds_increment_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] dds_increment_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // dds_increment_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> dds_increment_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          dds_increment_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // dds_increment_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> dds_increment_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          dds_increment_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                  // dds_increment_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> dds_increment_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] dds_increment_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                   // dds_increment_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> dds_increment_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          dds_increment_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                  // dds_increment_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> dds_increment_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                        // cpu_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid;                              // cpu_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                      // cpu_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [113:0] cpu_data_master_translator_avalon_universal_master_0_agent_cp_data;                               // cpu_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready;                              // addr_router:sink_ready -> cpu_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          vga_to_sdram_translator_avalon_universal_master_0_agent_cp_endofpacket;                           // vga_to_sdram_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          vga_to_sdram_translator_avalon_universal_master_0_agent_cp_valid;                                 // vga_to_sdram_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          vga_to_sdram_translator_avalon_universal_master_0_agent_cp_startofpacket;                         // vga_to_sdram_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [113:0] vga_to_sdram_translator_avalon_universal_master_0_agent_cp_data;                                  // vga_to_sdram_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          vga_to_sdram_translator_avalon_universal_master_0_agent_cp_ready;                                 // addr_router_001:sink_ready -> vga_to_sdram_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                 // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                       // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;               // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire  [113:0] cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                        // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                       // addr_router_002:sink_ready -> cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          addr_router_002_src_endofpacket;                                                                  // addr_router_002:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire          addr_router_002_src_valid;                                                                        // addr_router_002:src_valid -> limiter:cmd_sink_valid
	wire          addr_router_002_src_startofpacket;                                                                // addr_router_002:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [113:0] addr_router_002_src_data;                                                                         // addr_router_002:src_data -> limiter:cmd_sink_data
	wire   [24:0] addr_router_002_src_channel;                                                                      // addr_router_002:src_channel -> limiter:cmd_sink_channel
	wire          addr_router_002_src_ready;                                                                        // limiter:cmd_sink_ready -> addr_router_002:src_ready
	wire          limiter_rsp_src_endofpacket;                                                                      // limiter:rsp_src_endofpacket -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_rsp_src_valid;                                                                            // limiter:rsp_src_valid -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_rsp_src_startofpacket;                                                                    // limiter:rsp_src_startofpacket -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [113:0] limiter_rsp_src_data;                                                                             // limiter:rsp_src_data -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [24:0] limiter_rsp_src_channel;                                                                          // limiter:rsp_src_channel -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_rsp_src_ready;                                                                            // cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire          rst_controller_reset_out_reset;                                                                   // rst_controller:reset_out -> [agent_pipeline:reset, agent_pipeline_001:reset, agent_pipeline_002:reset, agent_pipeline_003:reset, agent_pipeline_004:reset, agent_pipeline_005:reset, agent_pipeline_006:reset, agent_pipeline_007:reset, agent_pipeline_008:reset, agent_pipeline_009:reset, agent_pipeline_010:reset, agent_pipeline_011:reset, agent_pipeline_014:reset, agent_pipeline_015:reset, agent_pipeline_016:reset, agent_pipeline_017:reset, agent_pipeline_018:reset, agent_pipeline_019:reset, agent_pipeline_020:reset, agent_pipeline_021:reset, agent_pipeline_022:reset, agent_pipeline_023:reset, agent_pipeline_024:reset, agent_pipeline_025:reset, agent_pipeline_026:reset, agent_pipeline_027:reset, agent_pipeline_032:reset, agent_pipeline_033:reset, agent_pipeline_034:reset, agent_pipeline_035:reset, agent_pipeline_038:reset, agent_pipeline_039:reset, agent_pipeline_040:reset, agent_pipeline_041:reset, agent_pipeline_044:reset, agent_pipeline_045:reset, agent_pipeline_046:reset, agent_pipeline_047:reset, agent_pipeline_048:reset, agent_pipeline_049:reset, audio:reset_reset_n, audio_data_fregen_s1_translator:reset, audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:reset, audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, audio_empty_s1_translator:reset, audio_empty_s1_translator_avalon_universal_slave_0_agent:reset, audio_empty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, audio_empty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, audio_fifo_full_s1_translator:reset, audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:reset, audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, audio_fifo_used_s1_translator:reset, audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:reset, audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, audio_out_data_audio_s1_translator:reset, audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:reset, audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, audio_out_pause_s1_translator:reset, audio_out_pause_s1_translator_avalon_universal_slave_0_agent:reset, audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, audio_out_stop_s1_translator:reset, audio_out_stop_s1_translator_avalon_universal_slave_0_agent:reset, audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, audio_sel:reset_n, audio_sel_s1_translator:reset, audio_sel_s1_translator_avalon_universal_slave_0_agent:reset, audio_sel_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, audio_sel_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, audio_wrclk_s1_translator:reset, audio_wrclk_s1_translator_avalon_universal_slave_0_agent:reset, audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, audio_wrreq_s1_translator:reset, audio_wrreq_s1_translator_avalon_universal_slave_0_agent:reset, audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, dds_increment:reset_n, dds_increment_s1_translator:reset, dds_increment_s1_translator_avalon_universal_slave_0_agent:reset, dds_increment_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, dds_increment_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, div_freq:reset_n, div_freq_s1_translator:reset, div_freq_s1_translator_avalon_universal_slave_0_agent:reset, div_freq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, div_freq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, id_router_016:reset, id_router_017:reset, id_router_019:reset, id_router_020:reset, id_router_022:reset, id_router_023:reset, id_router_024:reset, jtag_uart:rst_n, jtag_uart_avalon_jtag_slave_translator:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, key:reset_n, key_s1_translator:reset, key_s1_translator_avalon_universal_slave_0_agent:reset, key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, lfsr_clk_interrupt_gen:reset_n, lfsr_clk_interrupt_gen_s1_translator:reset, lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:reset, lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, lfsr_val:reset_n, lfsr_val_s1_translator:reset, lfsr_val_s1_translator_avalon_universal_slave_0_agent:reset, lfsr_val_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, lfsr_val_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, modulation_selector:reset_n, modulation_selector_s1_translator:reset, modulation_selector_s1_translator_avalon_universal_slave_0_agent:reset, modulation_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, modulation_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_016:reset, rsp_xbar_demux_017:reset, rsp_xbar_demux_019:reset, rsp_xbar_demux_020:reset, rsp_xbar_demux_022:reset, rsp_xbar_demux_023:reset, rsp_xbar_demux_024:reset, signal_selector:reset_n, signal_selector_s1_translator:reset, signal_selector_s1_translator_avalon_universal_slave_0_agent:reset, signal_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, signal_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sysid_qsys:reset_n, sysid_qsys_control_slave_translator:reset, sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer:reset_n, timer_s1_translator:reset, timer_s1_translator_avalon_universal_slave_0_agent:reset, timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire          rst_controller_001_reset_out_reset;                                                               // rst_controller_001:reset_out -> [addr_router:reset, addr_router_002:reset, agent_pipeline_012:reset, agent_pipeline_013:reset, cmd_xbar_demux:reset, cmd_xbar_demux_002:reset, cmd_xbar_mux_006:reset, cpu:reset_n, cpu_data_master_translator:reset, cpu_data_master_translator_avalon_universal_master_0_agent:reset, cpu_instruction_master_translator:reset, cpu_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu_jtag_debug_module_translator:reset, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, crosser:in_reset, crosser_001:in_reset, crosser_002:in_reset, crosser_003:in_reset, crosser_004:in_reset, crosser_005:out_reset, crosser_006:out_reset, crosser_007:out_reset, crosser_008:out_reset, crosser_009:out_reset, id_router_006:reset, irq_mapper:reset, irq_synchronizer:sender_reset, limiter:reset, limiter_pipeline:reset, limiter_pipeline_001:reset, rsp_xbar_demux_006:reset, rsp_xbar_mux:reset, rsp_xbar_mux_002:reset]
	wire          cpu_jtag_debug_module_reset_reset;                                                                // cpu:jtag_debug_module_resetrequest -> rst_controller_001:reset_in1
	wire          rst_controller_002_reset_out_reset;                                                               // rst_controller_002:reset_out -> [agent_pipeline_028:reset, agent_pipeline_029:reset, crosser:out_reset, crosser_005:in_reset, id_router_014:reset, keyboard_keys:reset_n, keyboard_keys_s1_translator:reset, keyboard_keys_s1_translator_avalon_universal_slave_0_agent:reset, keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_014:reset]
	wire          rst_controller_003_reset_out_reset;                                                               // rst_controller_003:reset_out -> [agent_pipeline_030:reset, agent_pipeline_031:reset, crosser_001:out_reset, crosser_006:in_reset, id_router_015:reset, mouse_pos:reset_n, mouse_pos_s1_translator:reset, mouse_pos_s1_translator_avalon_universal_slave_0_agent:reset, mouse_pos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, mouse_pos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_015:reset]
	wire          rst_controller_004_reset_out_reset;                                                               // rst_controller_004:reset_out -> [addr_router_001:reset, agent_pipeline_036:reset, agent_pipeline_037:reset, agent_pipeline_042:reset, agent_pipeline_043:reset, burst_adapter:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux_021:reset, crosser_002:out_reset, crosser_003:out_reset, crosser_004:out_reset, crosser_007:in_reset, crosser_008:in_reset, crosser_009:in_reset, id_router_018:reset, id_router_021:reset, rsp_xbar_demux_018:reset, rsp_xbar_demux_021:reset, sdram:reset_n, sdram_s1_translator:reset, sdram_s1_translator_avalon_universal_slave_0_agent:reset, sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, vga_to_nios_2_datamaster_translator:reset, vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:reset, vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, vga_to_sdram_translator:reset, vga_to_sdram_translator_avalon_universal_master_0_agent:reset, width_adapter:reset, width_adapter_001:reset]
	wire          cmd_xbar_demux_src0_endofpacket;                                                                  // cmd_xbar_demux:src0_endofpacket -> agent_pipeline:in_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                        // cmd_xbar_demux:src0_valid -> agent_pipeline:in_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                // cmd_xbar_demux:src0_startofpacket -> agent_pipeline:in_startofpacket
	wire  [113:0] cmd_xbar_demux_src0_data;                                                                         // cmd_xbar_demux:src0_data -> agent_pipeline:in_data
	wire   [24:0] cmd_xbar_demux_src0_channel;                                                                      // cmd_xbar_demux:src0_channel -> agent_pipeline:in_channel
	wire          cmd_xbar_demux_src1_endofpacket;                                                                  // cmd_xbar_demux:src1_endofpacket -> agent_pipeline_002:in_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                        // cmd_xbar_demux:src1_valid -> agent_pipeline_002:in_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                // cmd_xbar_demux:src1_startofpacket -> agent_pipeline_002:in_startofpacket
	wire  [113:0] cmd_xbar_demux_src1_data;                                                                         // cmd_xbar_demux:src1_data -> agent_pipeline_002:in_data
	wire   [24:0] cmd_xbar_demux_src1_channel;                                                                      // cmd_xbar_demux:src1_channel -> agent_pipeline_002:in_channel
	wire          cmd_xbar_demux_src2_endofpacket;                                                                  // cmd_xbar_demux:src2_endofpacket -> agent_pipeline_004:in_endofpacket
	wire          cmd_xbar_demux_src2_valid;                                                                        // cmd_xbar_demux:src2_valid -> agent_pipeline_004:in_valid
	wire          cmd_xbar_demux_src2_startofpacket;                                                                // cmd_xbar_demux:src2_startofpacket -> agent_pipeline_004:in_startofpacket
	wire  [113:0] cmd_xbar_demux_src2_data;                                                                         // cmd_xbar_demux:src2_data -> agent_pipeline_004:in_data
	wire   [24:0] cmd_xbar_demux_src2_channel;                                                                      // cmd_xbar_demux:src2_channel -> agent_pipeline_004:in_channel
	wire          cmd_xbar_demux_src3_endofpacket;                                                                  // cmd_xbar_demux:src3_endofpacket -> agent_pipeline_006:in_endofpacket
	wire          cmd_xbar_demux_src3_valid;                                                                        // cmd_xbar_demux:src3_valid -> agent_pipeline_006:in_valid
	wire          cmd_xbar_demux_src3_startofpacket;                                                                // cmd_xbar_demux:src3_startofpacket -> agent_pipeline_006:in_startofpacket
	wire  [113:0] cmd_xbar_demux_src3_data;                                                                         // cmd_xbar_demux:src3_data -> agent_pipeline_006:in_data
	wire   [24:0] cmd_xbar_demux_src3_channel;                                                                      // cmd_xbar_demux:src3_channel -> agent_pipeline_006:in_channel
	wire          cmd_xbar_demux_src4_endofpacket;                                                                  // cmd_xbar_demux:src4_endofpacket -> agent_pipeline_008:in_endofpacket
	wire          cmd_xbar_demux_src4_valid;                                                                        // cmd_xbar_demux:src4_valid -> agent_pipeline_008:in_valid
	wire          cmd_xbar_demux_src4_startofpacket;                                                                // cmd_xbar_demux:src4_startofpacket -> agent_pipeline_008:in_startofpacket
	wire  [113:0] cmd_xbar_demux_src4_data;                                                                         // cmd_xbar_demux:src4_data -> agent_pipeline_008:in_data
	wire   [24:0] cmd_xbar_demux_src4_channel;                                                                      // cmd_xbar_demux:src4_channel -> agent_pipeline_008:in_channel
	wire          cmd_xbar_demux_src5_endofpacket;                                                                  // cmd_xbar_demux:src5_endofpacket -> agent_pipeline_010:in_endofpacket
	wire          cmd_xbar_demux_src5_valid;                                                                        // cmd_xbar_demux:src5_valid -> agent_pipeline_010:in_valid
	wire          cmd_xbar_demux_src5_startofpacket;                                                                // cmd_xbar_demux:src5_startofpacket -> agent_pipeline_010:in_startofpacket
	wire  [113:0] cmd_xbar_demux_src5_data;                                                                         // cmd_xbar_demux:src5_data -> agent_pipeline_010:in_data
	wire   [24:0] cmd_xbar_demux_src5_channel;                                                                      // cmd_xbar_demux:src5_channel -> agent_pipeline_010:in_channel
	wire          cmd_xbar_demux_src6_endofpacket;                                                                  // cmd_xbar_demux:src6_endofpacket -> cmd_xbar_mux_006:sink0_endofpacket
	wire          cmd_xbar_demux_src6_valid;                                                                        // cmd_xbar_demux:src6_valid -> cmd_xbar_mux_006:sink0_valid
	wire          cmd_xbar_demux_src6_startofpacket;                                                                // cmd_xbar_demux:src6_startofpacket -> cmd_xbar_mux_006:sink0_startofpacket
	wire  [113:0] cmd_xbar_demux_src6_data;                                                                         // cmd_xbar_demux:src6_data -> cmd_xbar_mux_006:sink0_data
	wire   [24:0] cmd_xbar_demux_src6_channel;                                                                      // cmd_xbar_demux:src6_channel -> cmd_xbar_mux_006:sink0_channel
	wire          cmd_xbar_demux_src6_ready;                                                                        // cmd_xbar_mux_006:sink0_ready -> cmd_xbar_demux:src6_ready
	wire          cmd_xbar_demux_src7_endofpacket;                                                                  // cmd_xbar_demux:src7_endofpacket -> agent_pipeline_014:in_endofpacket
	wire          cmd_xbar_demux_src7_valid;                                                                        // cmd_xbar_demux:src7_valid -> agent_pipeline_014:in_valid
	wire          cmd_xbar_demux_src7_startofpacket;                                                                // cmd_xbar_demux:src7_startofpacket -> agent_pipeline_014:in_startofpacket
	wire  [113:0] cmd_xbar_demux_src7_data;                                                                         // cmd_xbar_demux:src7_data -> agent_pipeline_014:in_data
	wire   [24:0] cmd_xbar_demux_src7_channel;                                                                      // cmd_xbar_demux:src7_channel -> agent_pipeline_014:in_channel
	wire          cmd_xbar_demux_src8_endofpacket;                                                                  // cmd_xbar_demux:src8_endofpacket -> agent_pipeline_016:in_endofpacket
	wire          cmd_xbar_demux_src8_valid;                                                                        // cmd_xbar_demux:src8_valid -> agent_pipeline_016:in_valid
	wire          cmd_xbar_demux_src8_startofpacket;                                                                // cmd_xbar_demux:src8_startofpacket -> agent_pipeline_016:in_startofpacket
	wire  [113:0] cmd_xbar_demux_src8_data;                                                                         // cmd_xbar_demux:src8_data -> agent_pipeline_016:in_data
	wire   [24:0] cmd_xbar_demux_src8_channel;                                                                      // cmd_xbar_demux:src8_channel -> agent_pipeline_016:in_channel
	wire          cmd_xbar_demux_src9_endofpacket;                                                                  // cmd_xbar_demux:src9_endofpacket -> agent_pipeline_018:in_endofpacket
	wire          cmd_xbar_demux_src9_valid;                                                                        // cmd_xbar_demux:src9_valid -> agent_pipeline_018:in_valid
	wire          cmd_xbar_demux_src9_startofpacket;                                                                // cmd_xbar_demux:src9_startofpacket -> agent_pipeline_018:in_startofpacket
	wire  [113:0] cmd_xbar_demux_src9_data;                                                                         // cmd_xbar_demux:src9_data -> agent_pipeline_018:in_data
	wire   [24:0] cmd_xbar_demux_src9_channel;                                                                      // cmd_xbar_demux:src9_channel -> agent_pipeline_018:in_channel
	wire          cmd_xbar_demux_src10_endofpacket;                                                                 // cmd_xbar_demux:src10_endofpacket -> agent_pipeline_020:in_endofpacket
	wire          cmd_xbar_demux_src10_valid;                                                                       // cmd_xbar_demux:src10_valid -> agent_pipeline_020:in_valid
	wire          cmd_xbar_demux_src10_startofpacket;                                                               // cmd_xbar_demux:src10_startofpacket -> agent_pipeline_020:in_startofpacket
	wire  [113:0] cmd_xbar_demux_src10_data;                                                                        // cmd_xbar_demux:src10_data -> agent_pipeline_020:in_data
	wire   [24:0] cmd_xbar_demux_src10_channel;                                                                     // cmd_xbar_demux:src10_channel -> agent_pipeline_020:in_channel
	wire          cmd_xbar_demux_src11_endofpacket;                                                                 // cmd_xbar_demux:src11_endofpacket -> agent_pipeline_022:in_endofpacket
	wire          cmd_xbar_demux_src11_valid;                                                                       // cmd_xbar_demux:src11_valid -> agent_pipeline_022:in_valid
	wire          cmd_xbar_demux_src11_startofpacket;                                                               // cmd_xbar_demux:src11_startofpacket -> agent_pipeline_022:in_startofpacket
	wire  [113:0] cmd_xbar_demux_src11_data;                                                                        // cmd_xbar_demux:src11_data -> agent_pipeline_022:in_data
	wire   [24:0] cmd_xbar_demux_src11_channel;                                                                     // cmd_xbar_demux:src11_channel -> agent_pipeline_022:in_channel
	wire          cmd_xbar_demux_src12_endofpacket;                                                                 // cmd_xbar_demux:src12_endofpacket -> agent_pipeline_024:in_endofpacket
	wire          cmd_xbar_demux_src12_valid;                                                                       // cmd_xbar_demux:src12_valid -> agent_pipeline_024:in_valid
	wire          cmd_xbar_demux_src12_startofpacket;                                                               // cmd_xbar_demux:src12_startofpacket -> agent_pipeline_024:in_startofpacket
	wire  [113:0] cmd_xbar_demux_src12_data;                                                                        // cmd_xbar_demux:src12_data -> agent_pipeline_024:in_data
	wire   [24:0] cmd_xbar_demux_src12_channel;                                                                     // cmd_xbar_demux:src12_channel -> agent_pipeline_024:in_channel
	wire          cmd_xbar_demux_src13_endofpacket;                                                                 // cmd_xbar_demux:src13_endofpacket -> agent_pipeline_026:in_endofpacket
	wire          cmd_xbar_demux_src13_valid;                                                                       // cmd_xbar_demux:src13_valid -> agent_pipeline_026:in_valid
	wire          cmd_xbar_demux_src13_startofpacket;                                                               // cmd_xbar_demux:src13_startofpacket -> agent_pipeline_026:in_startofpacket
	wire  [113:0] cmd_xbar_demux_src13_data;                                                                        // cmd_xbar_demux:src13_data -> agent_pipeline_026:in_data
	wire   [24:0] cmd_xbar_demux_src13_channel;                                                                     // cmd_xbar_demux:src13_channel -> agent_pipeline_026:in_channel
	wire          cmd_xbar_demux_src16_endofpacket;                                                                 // cmd_xbar_demux:src16_endofpacket -> agent_pipeline_032:in_endofpacket
	wire          cmd_xbar_demux_src16_valid;                                                                       // cmd_xbar_demux:src16_valid -> agent_pipeline_032:in_valid
	wire          cmd_xbar_demux_src16_startofpacket;                                                               // cmd_xbar_demux:src16_startofpacket -> agent_pipeline_032:in_startofpacket
	wire  [113:0] cmd_xbar_demux_src16_data;                                                                        // cmd_xbar_demux:src16_data -> agent_pipeline_032:in_data
	wire   [24:0] cmd_xbar_demux_src16_channel;                                                                     // cmd_xbar_demux:src16_channel -> agent_pipeline_032:in_channel
	wire          cmd_xbar_demux_src17_endofpacket;                                                                 // cmd_xbar_demux:src17_endofpacket -> agent_pipeline_034:in_endofpacket
	wire          cmd_xbar_demux_src17_valid;                                                                       // cmd_xbar_demux:src17_valid -> agent_pipeline_034:in_valid
	wire          cmd_xbar_demux_src17_startofpacket;                                                               // cmd_xbar_demux:src17_startofpacket -> agent_pipeline_034:in_startofpacket
	wire  [113:0] cmd_xbar_demux_src17_data;                                                                        // cmd_xbar_demux:src17_data -> agent_pipeline_034:in_data
	wire   [24:0] cmd_xbar_demux_src17_channel;                                                                     // cmd_xbar_demux:src17_channel -> agent_pipeline_034:in_channel
	wire          cmd_xbar_demux_src19_endofpacket;                                                                 // cmd_xbar_demux:src19_endofpacket -> agent_pipeline_038:in_endofpacket
	wire          cmd_xbar_demux_src19_valid;                                                                       // cmd_xbar_demux:src19_valid -> agent_pipeline_038:in_valid
	wire          cmd_xbar_demux_src19_startofpacket;                                                               // cmd_xbar_demux:src19_startofpacket -> agent_pipeline_038:in_startofpacket
	wire  [113:0] cmd_xbar_demux_src19_data;                                                                        // cmd_xbar_demux:src19_data -> agent_pipeline_038:in_data
	wire   [24:0] cmd_xbar_demux_src19_channel;                                                                     // cmd_xbar_demux:src19_channel -> agent_pipeline_038:in_channel
	wire          cmd_xbar_demux_src20_endofpacket;                                                                 // cmd_xbar_demux:src20_endofpacket -> agent_pipeline_040:in_endofpacket
	wire          cmd_xbar_demux_src20_valid;                                                                       // cmd_xbar_demux:src20_valid -> agent_pipeline_040:in_valid
	wire          cmd_xbar_demux_src20_startofpacket;                                                               // cmd_xbar_demux:src20_startofpacket -> agent_pipeline_040:in_startofpacket
	wire  [113:0] cmd_xbar_demux_src20_data;                                                                        // cmd_xbar_demux:src20_data -> agent_pipeline_040:in_data
	wire   [24:0] cmd_xbar_demux_src20_channel;                                                                     // cmd_xbar_demux:src20_channel -> agent_pipeline_040:in_channel
	wire          cmd_xbar_demux_src22_endofpacket;                                                                 // cmd_xbar_demux:src22_endofpacket -> agent_pipeline_044:in_endofpacket
	wire          cmd_xbar_demux_src22_valid;                                                                       // cmd_xbar_demux:src22_valid -> agent_pipeline_044:in_valid
	wire          cmd_xbar_demux_src22_startofpacket;                                                               // cmd_xbar_demux:src22_startofpacket -> agent_pipeline_044:in_startofpacket
	wire  [113:0] cmd_xbar_demux_src22_data;                                                                        // cmd_xbar_demux:src22_data -> agent_pipeline_044:in_data
	wire   [24:0] cmd_xbar_demux_src22_channel;                                                                     // cmd_xbar_demux:src22_channel -> agent_pipeline_044:in_channel
	wire          cmd_xbar_demux_src23_endofpacket;                                                                 // cmd_xbar_demux:src23_endofpacket -> agent_pipeline_046:in_endofpacket
	wire          cmd_xbar_demux_src23_valid;                                                                       // cmd_xbar_demux:src23_valid -> agent_pipeline_046:in_valid
	wire          cmd_xbar_demux_src23_startofpacket;                                                               // cmd_xbar_demux:src23_startofpacket -> agent_pipeline_046:in_startofpacket
	wire  [113:0] cmd_xbar_demux_src23_data;                                                                        // cmd_xbar_demux:src23_data -> agent_pipeline_046:in_data
	wire   [24:0] cmd_xbar_demux_src23_channel;                                                                     // cmd_xbar_demux:src23_channel -> agent_pipeline_046:in_channel
	wire          cmd_xbar_demux_src24_endofpacket;                                                                 // cmd_xbar_demux:src24_endofpacket -> agent_pipeline_048:in_endofpacket
	wire          cmd_xbar_demux_src24_valid;                                                                       // cmd_xbar_demux:src24_valid -> agent_pipeline_048:in_valid
	wire          cmd_xbar_demux_src24_startofpacket;                                                               // cmd_xbar_demux:src24_startofpacket -> agent_pipeline_048:in_startofpacket
	wire  [113:0] cmd_xbar_demux_src24_data;                                                                        // cmd_xbar_demux:src24_data -> agent_pipeline_048:in_data
	wire   [24:0] cmd_xbar_demux_src24_channel;                                                                     // cmd_xbar_demux:src24_channel -> agent_pipeline_048:in_channel
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                              // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux_021:sink1_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                    // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux_021:sink1_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                            // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux_021:sink1_startofpacket
	wire  [113:0] cmd_xbar_demux_001_src0_data;                                                                     // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux_021:sink1_data
	wire   [24:0] cmd_xbar_demux_001_src0_channel;                                                                  // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux_021:sink1_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                    // cmd_xbar_mux_021:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_002_src0_endofpacket;                                                              // cmd_xbar_demux_002:src0_endofpacket -> cmd_xbar_mux_006:sink1_endofpacket
	wire          cmd_xbar_demux_002_src0_valid;                                                                    // cmd_xbar_demux_002:src0_valid -> cmd_xbar_mux_006:sink1_valid
	wire          cmd_xbar_demux_002_src0_startofpacket;                                                            // cmd_xbar_demux_002:src0_startofpacket -> cmd_xbar_mux_006:sink1_startofpacket
	wire  [113:0] cmd_xbar_demux_002_src0_data;                                                                     // cmd_xbar_demux_002:src0_data -> cmd_xbar_mux_006:sink1_data
	wire   [24:0] cmd_xbar_demux_002_src0_channel;                                                                  // cmd_xbar_demux_002:src0_channel -> cmd_xbar_mux_006:sink1_channel
	wire          cmd_xbar_demux_002_src0_ready;                                                                    // cmd_xbar_mux_006:sink1_ready -> cmd_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_src0_endofpacket;                                                                  // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                        // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [113:0] rsp_xbar_demux_src0_data;                                                                         // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [24:0] rsp_xbar_demux_src0_channel;                                                                      // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                        // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                              // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                    // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                            // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [113:0] rsp_xbar_demux_001_src0_data;                                                                     // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [24:0] rsp_xbar_demux_001_src0_channel;                                                                  // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                    // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                              // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                    // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                            // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [113:0] rsp_xbar_demux_002_src0_data;                                                                     // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire   [24:0] rsp_xbar_demux_002_src0_channel;                                                                  // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                    // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                              // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                    // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                            // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire  [113:0] rsp_xbar_demux_003_src0_data;                                                                     // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	wire   [24:0] rsp_xbar_demux_003_src0_channel;                                                                  // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                    // rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                              // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux:sink4_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                    // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux:sink4_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                            // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux:sink4_startofpacket
	wire  [113:0] rsp_xbar_demux_004_src0_data;                                                                     // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux:sink4_data
	wire   [24:0] rsp_xbar_demux_004_src0_channel;                                                                  // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux:sink4_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                    // rsp_xbar_mux:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                              // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux:sink5_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                    // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux:sink5_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                            // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux:sink5_startofpacket
	wire  [113:0] rsp_xbar_demux_005_src0_data;                                                                     // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux:sink5_data
	wire   [24:0] rsp_xbar_demux_005_src0_channel;                                                                  // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux:sink5_channel
	wire          rsp_xbar_demux_005_src0_ready;                                                                    // rsp_xbar_mux:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire          rsp_xbar_demux_006_src0_endofpacket;                                                              // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux:sink6_endofpacket
	wire          rsp_xbar_demux_006_src0_valid;                                                                    // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux:sink6_valid
	wire          rsp_xbar_demux_006_src0_startofpacket;                                                            // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux:sink6_startofpacket
	wire  [113:0] rsp_xbar_demux_006_src0_data;                                                                     // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux:sink6_data
	wire   [24:0] rsp_xbar_demux_006_src0_channel;                                                                  // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux:sink6_channel
	wire          rsp_xbar_demux_006_src0_ready;                                                                    // rsp_xbar_mux:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire          rsp_xbar_demux_006_src1_endofpacket;                                                              // rsp_xbar_demux_006:src1_endofpacket -> rsp_xbar_mux_002:sink0_endofpacket
	wire          rsp_xbar_demux_006_src1_valid;                                                                    // rsp_xbar_demux_006:src1_valid -> rsp_xbar_mux_002:sink0_valid
	wire          rsp_xbar_demux_006_src1_startofpacket;                                                            // rsp_xbar_demux_006:src1_startofpacket -> rsp_xbar_mux_002:sink0_startofpacket
	wire  [113:0] rsp_xbar_demux_006_src1_data;                                                                     // rsp_xbar_demux_006:src1_data -> rsp_xbar_mux_002:sink0_data
	wire   [24:0] rsp_xbar_demux_006_src1_channel;                                                                  // rsp_xbar_demux_006:src1_channel -> rsp_xbar_mux_002:sink0_channel
	wire          rsp_xbar_demux_006_src1_ready;                                                                    // rsp_xbar_mux_002:sink0_ready -> rsp_xbar_demux_006:src1_ready
	wire          rsp_xbar_demux_007_src0_endofpacket;                                                              // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux:sink7_endofpacket
	wire          rsp_xbar_demux_007_src0_valid;                                                                    // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux:sink7_valid
	wire          rsp_xbar_demux_007_src0_startofpacket;                                                            // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux:sink7_startofpacket
	wire  [113:0] rsp_xbar_demux_007_src0_data;                                                                     // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux:sink7_data
	wire   [24:0] rsp_xbar_demux_007_src0_channel;                                                                  // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux:sink7_channel
	wire          rsp_xbar_demux_007_src0_ready;                                                                    // rsp_xbar_mux:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire          rsp_xbar_demux_008_src0_endofpacket;                                                              // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux:sink8_endofpacket
	wire          rsp_xbar_demux_008_src0_valid;                                                                    // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux:sink8_valid
	wire          rsp_xbar_demux_008_src0_startofpacket;                                                            // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux:sink8_startofpacket
	wire  [113:0] rsp_xbar_demux_008_src0_data;                                                                     // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux:sink8_data
	wire   [24:0] rsp_xbar_demux_008_src0_channel;                                                                  // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux:sink8_channel
	wire          rsp_xbar_demux_008_src0_ready;                                                                    // rsp_xbar_mux:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire          rsp_xbar_demux_009_src0_endofpacket;                                                              // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux:sink9_endofpacket
	wire          rsp_xbar_demux_009_src0_valid;                                                                    // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux:sink9_valid
	wire          rsp_xbar_demux_009_src0_startofpacket;                                                            // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux:sink9_startofpacket
	wire  [113:0] rsp_xbar_demux_009_src0_data;                                                                     // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux:sink9_data
	wire   [24:0] rsp_xbar_demux_009_src0_channel;                                                                  // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux:sink9_channel
	wire          rsp_xbar_demux_009_src0_ready;                                                                    // rsp_xbar_mux:sink9_ready -> rsp_xbar_demux_009:src0_ready
	wire          rsp_xbar_demux_010_src0_endofpacket;                                                              // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux:sink10_endofpacket
	wire          rsp_xbar_demux_010_src0_valid;                                                                    // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux:sink10_valid
	wire          rsp_xbar_demux_010_src0_startofpacket;                                                            // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux:sink10_startofpacket
	wire  [113:0] rsp_xbar_demux_010_src0_data;                                                                     // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux:sink10_data
	wire   [24:0] rsp_xbar_demux_010_src0_channel;                                                                  // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux:sink10_channel
	wire          rsp_xbar_demux_010_src0_ready;                                                                    // rsp_xbar_mux:sink10_ready -> rsp_xbar_demux_010:src0_ready
	wire          rsp_xbar_demux_011_src0_endofpacket;                                                              // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux:sink11_endofpacket
	wire          rsp_xbar_demux_011_src0_valid;                                                                    // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux:sink11_valid
	wire          rsp_xbar_demux_011_src0_startofpacket;                                                            // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux:sink11_startofpacket
	wire  [113:0] rsp_xbar_demux_011_src0_data;                                                                     // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux:sink11_data
	wire   [24:0] rsp_xbar_demux_011_src0_channel;                                                                  // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux:sink11_channel
	wire          rsp_xbar_demux_011_src0_ready;                                                                    // rsp_xbar_mux:sink11_ready -> rsp_xbar_demux_011:src0_ready
	wire          rsp_xbar_demux_012_src0_endofpacket;                                                              // rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux:sink12_endofpacket
	wire          rsp_xbar_demux_012_src0_valid;                                                                    // rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux:sink12_valid
	wire          rsp_xbar_demux_012_src0_startofpacket;                                                            // rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux:sink12_startofpacket
	wire  [113:0] rsp_xbar_demux_012_src0_data;                                                                     // rsp_xbar_demux_012:src0_data -> rsp_xbar_mux:sink12_data
	wire   [24:0] rsp_xbar_demux_012_src0_channel;                                                                  // rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux:sink12_channel
	wire          rsp_xbar_demux_012_src0_ready;                                                                    // rsp_xbar_mux:sink12_ready -> rsp_xbar_demux_012:src0_ready
	wire          rsp_xbar_demux_013_src0_endofpacket;                                                              // rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux:sink13_endofpacket
	wire          rsp_xbar_demux_013_src0_valid;                                                                    // rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux:sink13_valid
	wire          rsp_xbar_demux_013_src0_startofpacket;                                                            // rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux:sink13_startofpacket
	wire  [113:0] rsp_xbar_demux_013_src0_data;                                                                     // rsp_xbar_demux_013:src0_data -> rsp_xbar_mux:sink13_data
	wire   [24:0] rsp_xbar_demux_013_src0_channel;                                                                  // rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux:sink13_channel
	wire          rsp_xbar_demux_013_src0_ready;                                                                    // rsp_xbar_mux:sink13_ready -> rsp_xbar_demux_013:src0_ready
	wire          rsp_xbar_demux_016_src0_endofpacket;                                                              // rsp_xbar_demux_016:src0_endofpacket -> rsp_xbar_mux:sink16_endofpacket
	wire          rsp_xbar_demux_016_src0_valid;                                                                    // rsp_xbar_demux_016:src0_valid -> rsp_xbar_mux:sink16_valid
	wire          rsp_xbar_demux_016_src0_startofpacket;                                                            // rsp_xbar_demux_016:src0_startofpacket -> rsp_xbar_mux:sink16_startofpacket
	wire  [113:0] rsp_xbar_demux_016_src0_data;                                                                     // rsp_xbar_demux_016:src0_data -> rsp_xbar_mux:sink16_data
	wire   [24:0] rsp_xbar_demux_016_src0_channel;                                                                  // rsp_xbar_demux_016:src0_channel -> rsp_xbar_mux:sink16_channel
	wire          rsp_xbar_demux_016_src0_ready;                                                                    // rsp_xbar_mux:sink16_ready -> rsp_xbar_demux_016:src0_ready
	wire          rsp_xbar_demux_017_src0_endofpacket;                                                              // rsp_xbar_demux_017:src0_endofpacket -> rsp_xbar_mux:sink17_endofpacket
	wire          rsp_xbar_demux_017_src0_valid;                                                                    // rsp_xbar_demux_017:src0_valid -> rsp_xbar_mux:sink17_valid
	wire          rsp_xbar_demux_017_src0_startofpacket;                                                            // rsp_xbar_demux_017:src0_startofpacket -> rsp_xbar_mux:sink17_startofpacket
	wire  [113:0] rsp_xbar_demux_017_src0_data;                                                                     // rsp_xbar_demux_017:src0_data -> rsp_xbar_mux:sink17_data
	wire   [24:0] rsp_xbar_demux_017_src0_channel;                                                                  // rsp_xbar_demux_017:src0_channel -> rsp_xbar_mux:sink17_channel
	wire          rsp_xbar_demux_017_src0_ready;                                                                    // rsp_xbar_mux:sink17_ready -> rsp_xbar_demux_017:src0_ready
	wire          rsp_xbar_demux_019_src0_endofpacket;                                                              // rsp_xbar_demux_019:src0_endofpacket -> rsp_xbar_mux:sink19_endofpacket
	wire          rsp_xbar_demux_019_src0_valid;                                                                    // rsp_xbar_demux_019:src0_valid -> rsp_xbar_mux:sink19_valid
	wire          rsp_xbar_demux_019_src0_startofpacket;                                                            // rsp_xbar_demux_019:src0_startofpacket -> rsp_xbar_mux:sink19_startofpacket
	wire  [113:0] rsp_xbar_demux_019_src0_data;                                                                     // rsp_xbar_demux_019:src0_data -> rsp_xbar_mux:sink19_data
	wire   [24:0] rsp_xbar_demux_019_src0_channel;                                                                  // rsp_xbar_demux_019:src0_channel -> rsp_xbar_mux:sink19_channel
	wire          rsp_xbar_demux_019_src0_ready;                                                                    // rsp_xbar_mux:sink19_ready -> rsp_xbar_demux_019:src0_ready
	wire          rsp_xbar_demux_020_src0_endofpacket;                                                              // rsp_xbar_demux_020:src0_endofpacket -> rsp_xbar_mux:sink20_endofpacket
	wire          rsp_xbar_demux_020_src0_valid;                                                                    // rsp_xbar_demux_020:src0_valid -> rsp_xbar_mux:sink20_valid
	wire          rsp_xbar_demux_020_src0_startofpacket;                                                            // rsp_xbar_demux_020:src0_startofpacket -> rsp_xbar_mux:sink20_startofpacket
	wire  [113:0] rsp_xbar_demux_020_src0_data;                                                                     // rsp_xbar_demux_020:src0_data -> rsp_xbar_mux:sink20_data
	wire   [24:0] rsp_xbar_demux_020_src0_channel;                                                                  // rsp_xbar_demux_020:src0_channel -> rsp_xbar_mux:sink20_channel
	wire          rsp_xbar_demux_020_src0_ready;                                                                    // rsp_xbar_mux:sink20_ready -> rsp_xbar_demux_020:src0_ready
	wire          rsp_xbar_demux_021_src1_endofpacket;                                                              // rsp_xbar_demux_021:src1_endofpacket -> vga_to_sdram_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_021_src1_valid;                                                                    // rsp_xbar_demux_021:src1_valid -> vga_to_sdram_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_021_src1_startofpacket;                                                            // rsp_xbar_demux_021:src1_startofpacket -> vga_to_sdram_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [113:0] rsp_xbar_demux_021_src1_data;                                                                     // rsp_xbar_demux_021:src1_data -> vga_to_sdram_translator_avalon_universal_master_0_agent:rp_data
	wire   [24:0] rsp_xbar_demux_021_src1_channel;                                                                  // rsp_xbar_demux_021:src1_channel -> vga_to_sdram_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_022_src0_endofpacket;                                                              // rsp_xbar_demux_022:src0_endofpacket -> rsp_xbar_mux:sink22_endofpacket
	wire          rsp_xbar_demux_022_src0_valid;                                                                    // rsp_xbar_demux_022:src0_valid -> rsp_xbar_mux:sink22_valid
	wire          rsp_xbar_demux_022_src0_startofpacket;                                                            // rsp_xbar_demux_022:src0_startofpacket -> rsp_xbar_mux:sink22_startofpacket
	wire  [113:0] rsp_xbar_demux_022_src0_data;                                                                     // rsp_xbar_demux_022:src0_data -> rsp_xbar_mux:sink22_data
	wire   [24:0] rsp_xbar_demux_022_src0_channel;                                                                  // rsp_xbar_demux_022:src0_channel -> rsp_xbar_mux:sink22_channel
	wire          rsp_xbar_demux_022_src0_ready;                                                                    // rsp_xbar_mux:sink22_ready -> rsp_xbar_demux_022:src0_ready
	wire          rsp_xbar_demux_023_src0_endofpacket;                                                              // rsp_xbar_demux_023:src0_endofpacket -> rsp_xbar_mux:sink23_endofpacket
	wire          rsp_xbar_demux_023_src0_valid;                                                                    // rsp_xbar_demux_023:src0_valid -> rsp_xbar_mux:sink23_valid
	wire          rsp_xbar_demux_023_src0_startofpacket;                                                            // rsp_xbar_demux_023:src0_startofpacket -> rsp_xbar_mux:sink23_startofpacket
	wire  [113:0] rsp_xbar_demux_023_src0_data;                                                                     // rsp_xbar_demux_023:src0_data -> rsp_xbar_mux:sink23_data
	wire   [24:0] rsp_xbar_demux_023_src0_channel;                                                                  // rsp_xbar_demux_023:src0_channel -> rsp_xbar_mux:sink23_channel
	wire          rsp_xbar_demux_023_src0_ready;                                                                    // rsp_xbar_mux:sink23_ready -> rsp_xbar_demux_023:src0_ready
	wire          rsp_xbar_demux_024_src0_endofpacket;                                                              // rsp_xbar_demux_024:src0_endofpacket -> rsp_xbar_mux:sink24_endofpacket
	wire          rsp_xbar_demux_024_src0_valid;                                                                    // rsp_xbar_demux_024:src0_valid -> rsp_xbar_mux:sink24_valid
	wire          rsp_xbar_demux_024_src0_startofpacket;                                                            // rsp_xbar_demux_024:src0_startofpacket -> rsp_xbar_mux:sink24_startofpacket
	wire  [113:0] rsp_xbar_demux_024_src0_data;                                                                     // rsp_xbar_demux_024:src0_data -> rsp_xbar_mux:sink24_data
	wire   [24:0] rsp_xbar_demux_024_src0_channel;                                                                  // rsp_xbar_demux_024:src0_channel -> rsp_xbar_mux:sink24_channel
	wire          rsp_xbar_demux_024_src0_ready;                                                                    // rsp_xbar_mux:sink24_ready -> rsp_xbar_demux_024:src0_ready
	wire          addr_router_src_endofpacket;                                                                      // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          addr_router_src_valid;                                                                            // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire          addr_router_src_startofpacket;                                                                    // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [113:0] addr_router_src_data;                                                                             // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire   [24:0] addr_router_src_channel;                                                                          // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire          addr_router_src_ready;                                                                            // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                     // rsp_xbar_mux:src_endofpacket -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                           // rsp_xbar_mux:src_valid -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                   // rsp_xbar_mux:src_startofpacket -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [113:0] rsp_xbar_mux_src_data;                                                                            // rsp_xbar_mux:src_data -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [24:0] rsp_xbar_mux_src_channel;                                                                         // rsp_xbar_mux:src_channel -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_src_ready;                                                                           // cpu_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	wire          addr_router_001_src_endofpacket;                                                                  // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          addr_router_001_src_valid;                                                                        // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire          addr_router_001_src_startofpacket;                                                                // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [113:0] addr_router_001_src_data;                                                                         // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire   [24:0] addr_router_001_src_channel;                                                                      // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire          addr_router_001_src_ready;                                                                        // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire          rsp_xbar_demux_021_src1_ready;                                                                    // vga_to_sdram_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_021:src1_ready
	wire          id_router_src_endofpacket;                                                                        // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                              // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                      // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [113:0] id_router_src_data;                                                                               // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [24:0] id_router_src_channel;                                                                            // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                              // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          id_router_001_src_endofpacket;                                                                    // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          id_router_001_src_valid;                                                                          // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire          id_router_001_src_startofpacket;                                                                  // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [113:0] id_router_001_src_data;                                                                           // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire   [24:0] id_router_001_src_channel;                                                                        // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire          id_router_001_src_ready;                                                                          // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire          id_router_002_src_endofpacket;                                                                    // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                          // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                                  // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [113:0] id_router_002_src_data;                                                                           // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire   [24:0] id_router_002_src_channel;                                                                        // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                          // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire          id_router_003_src_endofpacket;                                                                    // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                          // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                                  // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [113:0] id_router_003_src_data;                                                                           // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [24:0] id_router_003_src_channel;                                                                        // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                          // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          id_router_004_src_endofpacket;                                                                    // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          id_router_004_src_valid;                                                                          // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire          id_router_004_src_startofpacket;                                                                  // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [113:0] id_router_004_src_data;                                                                           // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire   [24:0] id_router_004_src_channel;                                                                        // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire          id_router_004_src_ready;                                                                          // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire          id_router_005_src_endofpacket;                                                                    // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          id_router_005_src_valid;                                                                          // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire          id_router_005_src_startofpacket;                                                                  // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [113:0] id_router_005_src_data;                                                                           // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [24:0] id_router_005_src_channel;                                                                        // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire          id_router_005_src_ready;                                                                          // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire          id_router_006_src_endofpacket;                                                                    // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire          id_router_006_src_valid;                                                                          // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire          id_router_006_src_startofpacket;                                                                  // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [113:0] id_router_006_src_data;                                                                           // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire   [24:0] id_router_006_src_channel;                                                                        // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire          id_router_006_src_ready;                                                                          // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire          id_router_007_src_endofpacket;                                                                    // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire          id_router_007_src_valid;                                                                          // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire          id_router_007_src_startofpacket;                                                                  // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [113:0] id_router_007_src_data;                                                                           // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire   [24:0] id_router_007_src_channel;                                                                        // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire          id_router_007_src_ready;                                                                          // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire          id_router_008_src_endofpacket;                                                                    // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire          id_router_008_src_valid;                                                                          // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire          id_router_008_src_startofpacket;                                                                  // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [113:0] id_router_008_src_data;                                                                           // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire   [24:0] id_router_008_src_channel;                                                                        // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire          id_router_008_src_ready;                                                                          // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire          id_router_009_src_endofpacket;                                                                    // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire          id_router_009_src_valid;                                                                          // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire          id_router_009_src_startofpacket;                                                                  // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [113:0] id_router_009_src_data;                                                                           // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire   [24:0] id_router_009_src_channel;                                                                        // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire          id_router_009_src_ready;                                                                          // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire          id_router_010_src_endofpacket;                                                                    // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire          id_router_010_src_valid;                                                                          // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire          id_router_010_src_startofpacket;                                                                  // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [113:0] id_router_010_src_data;                                                                           // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire   [24:0] id_router_010_src_channel;                                                                        // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire          id_router_010_src_ready;                                                                          // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire          id_router_011_src_endofpacket;                                                                    // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire          id_router_011_src_valid;                                                                          // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire          id_router_011_src_startofpacket;                                                                  // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire  [113:0] id_router_011_src_data;                                                                           // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire   [24:0] id_router_011_src_channel;                                                                        // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire          id_router_011_src_ready;                                                                          // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire          id_router_012_src_endofpacket;                                                                    // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire          id_router_012_src_valid;                                                                          // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire          id_router_012_src_startofpacket;                                                                  // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire  [113:0] id_router_012_src_data;                                                                           // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire   [24:0] id_router_012_src_channel;                                                                        // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire          id_router_012_src_ready;                                                                          // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire          id_router_013_src_endofpacket;                                                                    // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire          id_router_013_src_valid;                                                                          // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire          id_router_013_src_startofpacket;                                                                  // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire  [113:0] id_router_013_src_data;                                                                           // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire   [24:0] id_router_013_src_channel;                                                                        // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire          id_router_013_src_ready;                                                                          // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire          id_router_014_src_endofpacket;                                                                    // id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	wire          id_router_014_src_valid;                                                                          // id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	wire          id_router_014_src_startofpacket;                                                                  // id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	wire  [113:0] id_router_014_src_data;                                                                           // id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	wire   [24:0] id_router_014_src_channel;                                                                        // id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	wire          id_router_014_src_ready;                                                                          // rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	wire          id_router_015_src_endofpacket;                                                                    // id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	wire          id_router_015_src_valid;                                                                          // id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	wire          id_router_015_src_startofpacket;                                                                  // id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	wire  [113:0] id_router_015_src_data;                                                                           // id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	wire   [24:0] id_router_015_src_channel;                                                                        // id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	wire          id_router_015_src_ready;                                                                          // rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	wire          id_router_016_src_endofpacket;                                                                    // id_router_016:src_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	wire          id_router_016_src_valid;                                                                          // id_router_016:src_valid -> rsp_xbar_demux_016:sink_valid
	wire          id_router_016_src_startofpacket;                                                                  // id_router_016:src_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	wire  [113:0] id_router_016_src_data;                                                                           // id_router_016:src_data -> rsp_xbar_demux_016:sink_data
	wire   [24:0] id_router_016_src_channel;                                                                        // id_router_016:src_channel -> rsp_xbar_demux_016:sink_channel
	wire          id_router_016_src_ready;                                                                          // rsp_xbar_demux_016:sink_ready -> id_router_016:src_ready
	wire          id_router_017_src_endofpacket;                                                                    // id_router_017:src_endofpacket -> rsp_xbar_demux_017:sink_endofpacket
	wire          id_router_017_src_valid;                                                                          // id_router_017:src_valid -> rsp_xbar_demux_017:sink_valid
	wire          id_router_017_src_startofpacket;                                                                  // id_router_017:src_startofpacket -> rsp_xbar_demux_017:sink_startofpacket
	wire  [113:0] id_router_017_src_data;                                                                           // id_router_017:src_data -> rsp_xbar_demux_017:sink_data
	wire   [24:0] id_router_017_src_channel;                                                                        // id_router_017:src_channel -> rsp_xbar_demux_017:sink_channel
	wire          id_router_017_src_ready;                                                                          // rsp_xbar_demux_017:sink_ready -> id_router_017:src_ready
	wire          id_router_018_src_endofpacket;                                                                    // id_router_018:src_endofpacket -> rsp_xbar_demux_018:sink_endofpacket
	wire          id_router_018_src_valid;                                                                          // id_router_018:src_valid -> rsp_xbar_demux_018:sink_valid
	wire          id_router_018_src_startofpacket;                                                                  // id_router_018:src_startofpacket -> rsp_xbar_demux_018:sink_startofpacket
	wire  [113:0] id_router_018_src_data;                                                                           // id_router_018:src_data -> rsp_xbar_demux_018:sink_data
	wire   [24:0] id_router_018_src_channel;                                                                        // id_router_018:src_channel -> rsp_xbar_demux_018:sink_channel
	wire          id_router_018_src_ready;                                                                          // rsp_xbar_demux_018:sink_ready -> id_router_018:src_ready
	wire          id_router_019_src_endofpacket;                                                                    // id_router_019:src_endofpacket -> rsp_xbar_demux_019:sink_endofpacket
	wire          id_router_019_src_valid;                                                                          // id_router_019:src_valid -> rsp_xbar_demux_019:sink_valid
	wire          id_router_019_src_startofpacket;                                                                  // id_router_019:src_startofpacket -> rsp_xbar_demux_019:sink_startofpacket
	wire  [113:0] id_router_019_src_data;                                                                           // id_router_019:src_data -> rsp_xbar_demux_019:sink_data
	wire   [24:0] id_router_019_src_channel;                                                                        // id_router_019:src_channel -> rsp_xbar_demux_019:sink_channel
	wire          id_router_019_src_ready;                                                                          // rsp_xbar_demux_019:sink_ready -> id_router_019:src_ready
	wire          id_router_020_src_endofpacket;                                                                    // id_router_020:src_endofpacket -> rsp_xbar_demux_020:sink_endofpacket
	wire          id_router_020_src_valid;                                                                          // id_router_020:src_valid -> rsp_xbar_demux_020:sink_valid
	wire          id_router_020_src_startofpacket;                                                                  // id_router_020:src_startofpacket -> rsp_xbar_demux_020:sink_startofpacket
	wire  [113:0] id_router_020_src_data;                                                                           // id_router_020:src_data -> rsp_xbar_demux_020:sink_data
	wire   [24:0] id_router_020_src_channel;                                                                        // id_router_020:src_channel -> rsp_xbar_demux_020:sink_channel
	wire          id_router_020_src_ready;                                                                          // rsp_xbar_demux_020:sink_ready -> id_router_020:src_ready
	wire          id_router_022_src_endofpacket;                                                                    // id_router_022:src_endofpacket -> rsp_xbar_demux_022:sink_endofpacket
	wire          id_router_022_src_valid;                                                                          // id_router_022:src_valid -> rsp_xbar_demux_022:sink_valid
	wire          id_router_022_src_startofpacket;                                                                  // id_router_022:src_startofpacket -> rsp_xbar_demux_022:sink_startofpacket
	wire  [113:0] id_router_022_src_data;                                                                           // id_router_022:src_data -> rsp_xbar_demux_022:sink_data
	wire   [24:0] id_router_022_src_channel;                                                                        // id_router_022:src_channel -> rsp_xbar_demux_022:sink_channel
	wire          id_router_022_src_ready;                                                                          // rsp_xbar_demux_022:sink_ready -> id_router_022:src_ready
	wire          id_router_023_src_endofpacket;                                                                    // id_router_023:src_endofpacket -> rsp_xbar_demux_023:sink_endofpacket
	wire          id_router_023_src_valid;                                                                          // id_router_023:src_valid -> rsp_xbar_demux_023:sink_valid
	wire          id_router_023_src_startofpacket;                                                                  // id_router_023:src_startofpacket -> rsp_xbar_demux_023:sink_startofpacket
	wire  [113:0] id_router_023_src_data;                                                                           // id_router_023:src_data -> rsp_xbar_demux_023:sink_data
	wire   [24:0] id_router_023_src_channel;                                                                        // id_router_023:src_channel -> rsp_xbar_demux_023:sink_channel
	wire          id_router_023_src_ready;                                                                          // rsp_xbar_demux_023:sink_ready -> id_router_023:src_ready
	wire          id_router_024_src_endofpacket;                                                                    // id_router_024:src_endofpacket -> rsp_xbar_demux_024:sink_endofpacket
	wire          id_router_024_src_valid;                                                                          // id_router_024:src_valid -> rsp_xbar_demux_024:sink_valid
	wire          id_router_024_src_startofpacket;                                                                  // id_router_024:src_startofpacket -> rsp_xbar_demux_024:sink_startofpacket
	wire  [113:0] id_router_024_src_data;                                                                           // id_router_024:src_data -> rsp_xbar_demux_024:sink_data
	wire   [24:0] id_router_024_src_channel;                                                                        // id_router_024:src_channel -> rsp_xbar_demux_024:sink_channel
	wire          id_router_024_src_ready;                                                                          // rsp_xbar_demux_024:sink_ready -> id_router_024:src_ready
	wire          cmd_xbar_mux_021_src_endofpacket;                                                                 // cmd_xbar_mux_021:src_endofpacket -> width_adapter:in_endofpacket
	wire          cmd_xbar_mux_021_src_valid;                                                                       // cmd_xbar_mux_021:src_valid -> width_adapter:in_valid
	wire          cmd_xbar_mux_021_src_startofpacket;                                                               // cmd_xbar_mux_021:src_startofpacket -> width_adapter:in_startofpacket
	wire  [113:0] cmd_xbar_mux_021_src_data;                                                                        // cmd_xbar_mux_021:src_data -> width_adapter:in_data
	wire   [24:0] cmd_xbar_mux_021_src_channel;                                                                     // cmd_xbar_mux_021:src_channel -> width_adapter:in_channel
	wire          cmd_xbar_mux_021_src_ready;                                                                       // width_adapter:in_ready -> cmd_xbar_mux_021:src_ready
	wire          width_adapter_src_endofpacket;                                                                    // width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	wire          width_adapter_src_valid;                                                                          // width_adapter:out_valid -> burst_adapter:sink0_valid
	wire          width_adapter_src_startofpacket;                                                                  // width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	wire   [95:0] width_adapter_src_data;                                                                           // width_adapter:out_data -> burst_adapter:sink0_data
	wire          width_adapter_src_ready;                                                                          // burst_adapter:sink0_ready -> width_adapter:out_ready
	wire   [24:0] width_adapter_src_channel;                                                                        // width_adapter:out_channel -> burst_adapter:sink0_channel
	wire          id_router_021_src_endofpacket;                                                                    // id_router_021:src_endofpacket -> width_adapter_001:in_endofpacket
	wire          id_router_021_src_valid;                                                                          // id_router_021:src_valid -> width_adapter_001:in_valid
	wire          id_router_021_src_startofpacket;                                                                  // id_router_021:src_startofpacket -> width_adapter_001:in_startofpacket
	wire   [95:0] id_router_021_src_data;                                                                           // id_router_021:src_data -> width_adapter_001:in_data
	wire   [24:0] id_router_021_src_channel;                                                                        // id_router_021:src_channel -> width_adapter_001:in_channel
	wire          id_router_021_src_ready;                                                                          // width_adapter_001:in_ready -> id_router_021:src_ready
	wire          width_adapter_001_src_endofpacket;                                                                // width_adapter_001:out_endofpacket -> rsp_xbar_demux_021:sink_endofpacket
	wire          width_adapter_001_src_valid;                                                                      // width_adapter_001:out_valid -> rsp_xbar_demux_021:sink_valid
	wire          width_adapter_001_src_startofpacket;                                                              // width_adapter_001:out_startofpacket -> rsp_xbar_demux_021:sink_startofpacket
	wire  [113:0] width_adapter_001_src_data;                                                                       // width_adapter_001:out_data -> rsp_xbar_demux_021:sink_data
	wire          width_adapter_001_src_ready;                                                                      // rsp_xbar_demux_021:sink_ready -> width_adapter_001:out_ready
	wire   [24:0] width_adapter_001_src_channel;                                                                    // width_adapter_001:out_channel -> rsp_xbar_demux_021:sink_channel
	wire          crosser_out_endofpacket;                                                                          // crosser:out_endofpacket -> agent_pipeline_028:in_endofpacket
	wire          crosser_out_valid;                                                                                // crosser:out_valid -> agent_pipeline_028:in_valid
	wire          crosser_out_startofpacket;                                                                        // crosser:out_startofpacket -> agent_pipeline_028:in_startofpacket
	wire  [113:0] crosser_out_data;                                                                                 // crosser:out_data -> agent_pipeline_028:in_data
	wire   [24:0] crosser_out_channel;                                                                              // crosser:out_channel -> agent_pipeline_028:in_channel
	wire          cmd_xbar_demux_src14_endofpacket;                                                                 // cmd_xbar_demux:src14_endofpacket -> crosser:in_endofpacket
	wire          cmd_xbar_demux_src14_valid;                                                                       // cmd_xbar_demux:src14_valid -> crosser:in_valid
	wire          cmd_xbar_demux_src14_startofpacket;                                                               // cmd_xbar_demux:src14_startofpacket -> crosser:in_startofpacket
	wire  [113:0] cmd_xbar_demux_src14_data;                                                                        // cmd_xbar_demux:src14_data -> crosser:in_data
	wire   [24:0] cmd_xbar_demux_src14_channel;                                                                     // cmd_xbar_demux:src14_channel -> crosser:in_channel
	wire          cmd_xbar_demux_src14_ready;                                                                       // crosser:in_ready -> cmd_xbar_demux:src14_ready
	wire          crosser_001_out_endofpacket;                                                                      // crosser_001:out_endofpacket -> agent_pipeline_030:in_endofpacket
	wire          crosser_001_out_valid;                                                                            // crosser_001:out_valid -> agent_pipeline_030:in_valid
	wire          crosser_001_out_startofpacket;                                                                    // crosser_001:out_startofpacket -> agent_pipeline_030:in_startofpacket
	wire  [113:0] crosser_001_out_data;                                                                             // crosser_001:out_data -> agent_pipeline_030:in_data
	wire   [24:0] crosser_001_out_channel;                                                                          // crosser_001:out_channel -> agent_pipeline_030:in_channel
	wire          cmd_xbar_demux_src15_endofpacket;                                                                 // cmd_xbar_demux:src15_endofpacket -> crosser_001:in_endofpacket
	wire          cmd_xbar_demux_src15_valid;                                                                       // cmd_xbar_demux:src15_valid -> crosser_001:in_valid
	wire          cmd_xbar_demux_src15_startofpacket;                                                               // cmd_xbar_demux:src15_startofpacket -> crosser_001:in_startofpacket
	wire  [113:0] cmd_xbar_demux_src15_data;                                                                        // cmd_xbar_demux:src15_data -> crosser_001:in_data
	wire   [24:0] cmd_xbar_demux_src15_channel;                                                                     // cmd_xbar_demux:src15_channel -> crosser_001:in_channel
	wire          cmd_xbar_demux_src15_ready;                                                                       // crosser_001:in_ready -> cmd_xbar_demux:src15_ready
	wire          crosser_002_out_endofpacket;                                                                      // crosser_002:out_endofpacket -> agent_pipeline_036:in_endofpacket
	wire          crosser_002_out_valid;                                                                            // crosser_002:out_valid -> agent_pipeline_036:in_valid
	wire          crosser_002_out_startofpacket;                                                                    // crosser_002:out_startofpacket -> agent_pipeline_036:in_startofpacket
	wire  [113:0] crosser_002_out_data;                                                                             // crosser_002:out_data -> agent_pipeline_036:in_data
	wire   [24:0] crosser_002_out_channel;                                                                          // crosser_002:out_channel -> agent_pipeline_036:in_channel
	wire          cmd_xbar_demux_src18_endofpacket;                                                                 // cmd_xbar_demux:src18_endofpacket -> crosser_002:in_endofpacket
	wire          cmd_xbar_demux_src18_valid;                                                                       // cmd_xbar_demux:src18_valid -> crosser_002:in_valid
	wire          cmd_xbar_demux_src18_startofpacket;                                                               // cmd_xbar_demux:src18_startofpacket -> crosser_002:in_startofpacket
	wire  [113:0] cmd_xbar_demux_src18_data;                                                                        // cmd_xbar_demux:src18_data -> crosser_002:in_data
	wire   [24:0] cmd_xbar_demux_src18_channel;                                                                     // cmd_xbar_demux:src18_channel -> crosser_002:in_channel
	wire          cmd_xbar_demux_src18_ready;                                                                       // crosser_002:in_ready -> cmd_xbar_demux:src18_ready
	wire          crosser_003_out_endofpacket;                                                                      // crosser_003:out_endofpacket -> cmd_xbar_mux_021:sink0_endofpacket
	wire          crosser_003_out_valid;                                                                            // crosser_003:out_valid -> cmd_xbar_mux_021:sink0_valid
	wire          crosser_003_out_startofpacket;                                                                    // crosser_003:out_startofpacket -> cmd_xbar_mux_021:sink0_startofpacket
	wire  [113:0] crosser_003_out_data;                                                                             // crosser_003:out_data -> cmd_xbar_mux_021:sink0_data
	wire   [24:0] crosser_003_out_channel;                                                                          // crosser_003:out_channel -> cmd_xbar_mux_021:sink0_channel
	wire          crosser_003_out_ready;                                                                            // cmd_xbar_mux_021:sink0_ready -> crosser_003:out_ready
	wire          cmd_xbar_demux_src21_endofpacket;                                                                 // cmd_xbar_demux:src21_endofpacket -> crosser_003:in_endofpacket
	wire          cmd_xbar_demux_src21_valid;                                                                       // cmd_xbar_demux:src21_valid -> crosser_003:in_valid
	wire          cmd_xbar_demux_src21_startofpacket;                                                               // cmd_xbar_demux:src21_startofpacket -> crosser_003:in_startofpacket
	wire  [113:0] cmd_xbar_demux_src21_data;                                                                        // cmd_xbar_demux:src21_data -> crosser_003:in_data
	wire   [24:0] cmd_xbar_demux_src21_channel;                                                                     // cmd_xbar_demux:src21_channel -> crosser_003:in_channel
	wire          cmd_xbar_demux_src21_ready;                                                                       // crosser_003:in_ready -> cmd_xbar_demux:src21_ready
	wire          crosser_004_out_endofpacket;                                                                      // crosser_004:out_endofpacket -> cmd_xbar_mux_021:sink2_endofpacket
	wire          crosser_004_out_valid;                                                                            // crosser_004:out_valid -> cmd_xbar_mux_021:sink2_valid
	wire          crosser_004_out_startofpacket;                                                                    // crosser_004:out_startofpacket -> cmd_xbar_mux_021:sink2_startofpacket
	wire  [113:0] crosser_004_out_data;                                                                             // crosser_004:out_data -> cmd_xbar_mux_021:sink2_data
	wire   [24:0] crosser_004_out_channel;                                                                          // crosser_004:out_channel -> cmd_xbar_mux_021:sink2_channel
	wire          crosser_004_out_ready;                                                                            // cmd_xbar_mux_021:sink2_ready -> crosser_004:out_ready
	wire          cmd_xbar_demux_002_src1_endofpacket;                                                              // cmd_xbar_demux_002:src1_endofpacket -> crosser_004:in_endofpacket
	wire          cmd_xbar_demux_002_src1_valid;                                                                    // cmd_xbar_demux_002:src1_valid -> crosser_004:in_valid
	wire          cmd_xbar_demux_002_src1_startofpacket;                                                            // cmd_xbar_demux_002:src1_startofpacket -> crosser_004:in_startofpacket
	wire  [113:0] cmd_xbar_demux_002_src1_data;                                                                     // cmd_xbar_demux_002:src1_data -> crosser_004:in_data
	wire   [24:0] cmd_xbar_demux_002_src1_channel;                                                                  // cmd_xbar_demux_002:src1_channel -> crosser_004:in_channel
	wire          cmd_xbar_demux_002_src1_ready;                                                                    // crosser_004:in_ready -> cmd_xbar_demux_002:src1_ready
	wire          crosser_005_out_endofpacket;                                                                      // crosser_005:out_endofpacket -> rsp_xbar_mux:sink14_endofpacket
	wire          crosser_005_out_valid;                                                                            // crosser_005:out_valid -> rsp_xbar_mux:sink14_valid
	wire          crosser_005_out_startofpacket;                                                                    // crosser_005:out_startofpacket -> rsp_xbar_mux:sink14_startofpacket
	wire  [113:0] crosser_005_out_data;                                                                             // crosser_005:out_data -> rsp_xbar_mux:sink14_data
	wire   [24:0] crosser_005_out_channel;                                                                          // crosser_005:out_channel -> rsp_xbar_mux:sink14_channel
	wire          crosser_005_out_ready;                                                                            // rsp_xbar_mux:sink14_ready -> crosser_005:out_ready
	wire          rsp_xbar_demux_014_src0_endofpacket;                                                              // rsp_xbar_demux_014:src0_endofpacket -> crosser_005:in_endofpacket
	wire          rsp_xbar_demux_014_src0_valid;                                                                    // rsp_xbar_demux_014:src0_valid -> crosser_005:in_valid
	wire          rsp_xbar_demux_014_src0_startofpacket;                                                            // rsp_xbar_demux_014:src0_startofpacket -> crosser_005:in_startofpacket
	wire  [113:0] rsp_xbar_demux_014_src0_data;                                                                     // rsp_xbar_demux_014:src0_data -> crosser_005:in_data
	wire   [24:0] rsp_xbar_demux_014_src0_channel;                                                                  // rsp_xbar_demux_014:src0_channel -> crosser_005:in_channel
	wire          rsp_xbar_demux_014_src0_ready;                                                                    // crosser_005:in_ready -> rsp_xbar_demux_014:src0_ready
	wire          crosser_006_out_endofpacket;                                                                      // crosser_006:out_endofpacket -> rsp_xbar_mux:sink15_endofpacket
	wire          crosser_006_out_valid;                                                                            // crosser_006:out_valid -> rsp_xbar_mux:sink15_valid
	wire          crosser_006_out_startofpacket;                                                                    // crosser_006:out_startofpacket -> rsp_xbar_mux:sink15_startofpacket
	wire  [113:0] crosser_006_out_data;                                                                             // crosser_006:out_data -> rsp_xbar_mux:sink15_data
	wire   [24:0] crosser_006_out_channel;                                                                          // crosser_006:out_channel -> rsp_xbar_mux:sink15_channel
	wire          crosser_006_out_ready;                                                                            // rsp_xbar_mux:sink15_ready -> crosser_006:out_ready
	wire          rsp_xbar_demux_015_src0_endofpacket;                                                              // rsp_xbar_demux_015:src0_endofpacket -> crosser_006:in_endofpacket
	wire          rsp_xbar_demux_015_src0_valid;                                                                    // rsp_xbar_demux_015:src0_valid -> crosser_006:in_valid
	wire          rsp_xbar_demux_015_src0_startofpacket;                                                            // rsp_xbar_demux_015:src0_startofpacket -> crosser_006:in_startofpacket
	wire  [113:0] rsp_xbar_demux_015_src0_data;                                                                     // rsp_xbar_demux_015:src0_data -> crosser_006:in_data
	wire   [24:0] rsp_xbar_demux_015_src0_channel;                                                                  // rsp_xbar_demux_015:src0_channel -> crosser_006:in_channel
	wire          rsp_xbar_demux_015_src0_ready;                                                                    // crosser_006:in_ready -> rsp_xbar_demux_015:src0_ready
	wire          crosser_007_out_endofpacket;                                                                      // crosser_007:out_endofpacket -> rsp_xbar_mux:sink18_endofpacket
	wire          crosser_007_out_valid;                                                                            // crosser_007:out_valid -> rsp_xbar_mux:sink18_valid
	wire          crosser_007_out_startofpacket;                                                                    // crosser_007:out_startofpacket -> rsp_xbar_mux:sink18_startofpacket
	wire  [113:0] crosser_007_out_data;                                                                             // crosser_007:out_data -> rsp_xbar_mux:sink18_data
	wire   [24:0] crosser_007_out_channel;                                                                          // crosser_007:out_channel -> rsp_xbar_mux:sink18_channel
	wire          crosser_007_out_ready;                                                                            // rsp_xbar_mux:sink18_ready -> crosser_007:out_ready
	wire          rsp_xbar_demux_018_src0_endofpacket;                                                              // rsp_xbar_demux_018:src0_endofpacket -> crosser_007:in_endofpacket
	wire          rsp_xbar_demux_018_src0_valid;                                                                    // rsp_xbar_demux_018:src0_valid -> crosser_007:in_valid
	wire          rsp_xbar_demux_018_src0_startofpacket;                                                            // rsp_xbar_demux_018:src0_startofpacket -> crosser_007:in_startofpacket
	wire  [113:0] rsp_xbar_demux_018_src0_data;                                                                     // rsp_xbar_demux_018:src0_data -> crosser_007:in_data
	wire   [24:0] rsp_xbar_demux_018_src0_channel;                                                                  // rsp_xbar_demux_018:src0_channel -> crosser_007:in_channel
	wire          rsp_xbar_demux_018_src0_ready;                                                                    // crosser_007:in_ready -> rsp_xbar_demux_018:src0_ready
	wire          crosser_008_out_endofpacket;                                                                      // crosser_008:out_endofpacket -> rsp_xbar_mux:sink21_endofpacket
	wire          crosser_008_out_valid;                                                                            // crosser_008:out_valid -> rsp_xbar_mux:sink21_valid
	wire          crosser_008_out_startofpacket;                                                                    // crosser_008:out_startofpacket -> rsp_xbar_mux:sink21_startofpacket
	wire  [113:0] crosser_008_out_data;                                                                             // crosser_008:out_data -> rsp_xbar_mux:sink21_data
	wire   [24:0] crosser_008_out_channel;                                                                          // crosser_008:out_channel -> rsp_xbar_mux:sink21_channel
	wire          crosser_008_out_ready;                                                                            // rsp_xbar_mux:sink21_ready -> crosser_008:out_ready
	wire          rsp_xbar_demux_021_src0_endofpacket;                                                              // rsp_xbar_demux_021:src0_endofpacket -> crosser_008:in_endofpacket
	wire          rsp_xbar_demux_021_src0_valid;                                                                    // rsp_xbar_demux_021:src0_valid -> crosser_008:in_valid
	wire          rsp_xbar_demux_021_src0_startofpacket;                                                            // rsp_xbar_demux_021:src0_startofpacket -> crosser_008:in_startofpacket
	wire  [113:0] rsp_xbar_demux_021_src0_data;                                                                     // rsp_xbar_demux_021:src0_data -> crosser_008:in_data
	wire   [24:0] rsp_xbar_demux_021_src0_channel;                                                                  // rsp_xbar_demux_021:src0_channel -> crosser_008:in_channel
	wire          rsp_xbar_demux_021_src0_ready;                                                                    // crosser_008:in_ready -> rsp_xbar_demux_021:src0_ready
	wire          crosser_009_out_endofpacket;                                                                      // crosser_009:out_endofpacket -> rsp_xbar_mux_002:sink1_endofpacket
	wire          crosser_009_out_valid;                                                                            // crosser_009:out_valid -> rsp_xbar_mux_002:sink1_valid
	wire          crosser_009_out_startofpacket;                                                                    // crosser_009:out_startofpacket -> rsp_xbar_mux_002:sink1_startofpacket
	wire  [113:0] crosser_009_out_data;                                                                             // crosser_009:out_data -> rsp_xbar_mux_002:sink1_data
	wire   [24:0] crosser_009_out_channel;                                                                          // crosser_009:out_channel -> rsp_xbar_mux_002:sink1_channel
	wire          crosser_009_out_ready;                                                                            // rsp_xbar_mux_002:sink1_ready -> crosser_009:out_ready
	wire          rsp_xbar_demux_021_src2_endofpacket;                                                              // rsp_xbar_demux_021:src2_endofpacket -> crosser_009:in_endofpacket
	wire          rsp_xbar_demux_021_src2_valid;                                                                    // rsp_xbar_demux_021:src2_valid -> crosser_009:in_valid
	wire          rsp_xbar_demux_021_src2_startofpacket;                                                            // rsp_xbar_demux_021:src2_startofpacket -> crosser_009:in_startofpacket
	wire  [113:0] rsp_xbar_demux_021_src2_data;                                                                     // rsp_xbar_demux_021:src2_data -> crosser_009:in_data
	wire   [24:0] rsp_xbar_demux_021_src2_channel;                                                                  // rsp_xbar_demux_021:src2_channel -> crosser_009:in_channel
	wire          rsp_xbar_demux_021_src2_ready;                                                                    // crosser_009:in_ready -> rsp_xbar_demux_021:src2_ready
	wire          limiter_pipeline_source0_endofpacket;                                                             // limiter_pipeline:out_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire          limiter_pipeline_source0_valid;                                                                   // limiter_pipeline:out_valid -> cmd_xbar_demux_002:sink_valid
	wire          limiter_pipeline_source0_startofpacket;                                                           // limiter_pipeline:out_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire  [113:0] limiter_pipeline_source0_data;                                                                    // limiter_pipeline:out_data -> cmd_xbar_demux_002:sink_data
	wire   [24:0] limiter_pipeline_source0_channel;                                                                 // limiter_pipeline:out_channel -> cmd_xbar_demux_002:sink_channel
	wire          limiter_pipeline_source0_ready;                                                                   // cmd_xbar_demux_002:sink_ready -> limiter_pipeline:out_ready
	wire          limiter_cmd_src_endofpacket;                                                                      // limiter:cmd_src_endofpacket -> limiter_pipeline:in_endofpacket
	wire    [0:0] limiter_cmd_src_valid;                                                                            // limiter:cmd_src_valid -> limiter_pipeline:in_valid
	wire          limiter_cmd_src_startofpacket;                                                                    // limiter:cmd_src_startofpacket -> limiter_pipeline:in_startofpacket
	wire  [113:0] limiter_cmd_src_data;                                                                             // limiter:cmd_src_data -> limiter_pipeline:in_data
	wire   [24:0] limiter_cmd_src_channel;                                                                          // limiter:cmd_src_channel -> limiter_pipeline:in_channel
	wire          limiter_cmd_src_ready;                                                                            // limiter_pipeline:in_ready -> limiter:cmd_src_ready
	wire          rsp_xbar_mux_002_src_endofpacket;                                                                 // rsp_xbar_mux_002:src_endofpacket -> limiter_pipeline_001:in_endofpacket
	wire          rsp_xbar_mux_002_src_valid;                                                                       // rsp_xbar_mux_002:src_valid -> limiter_pipeline_001:in_valid
	wire          rsp_xbar_mux_002_src_startofpacket;                                                               // rsp_xbar_mux_002:src_startofpacket -> limiter_pipeline_001:in_startofpacket
	wire  [113:0] rsp_xbar_mux_002_src_data;                                                                        // rsp_xbar_mux_002:src_data -> limiter_pipeline_001:in_data
	wire   [24:0] rsp_xbar_mux_002_src_channel;                                                                     // rsp_xbar_mux_002:src_channel -> limiter_pipeline_001:in_channel
	wire          rsp_xbar_mux_002_src_ready;                                                                       // limiter_pipeline_001:in_ready -> rsp_xbar_mux_002:src_ready
	wire          limiter_pipeline_001_source0_endofpacket;                                                         // limiter_pipeline_001:out_endofpacket -> limiter:rsp_sink_endofpacket
	wire          limiter_pipeline_001_source0_valid;                                                               // limiter_pipeline_001:out_valid -> limiter:rsp_sink_valid
	wire          limiter_pipeline_001_source0_startofpacket;                                                       // limiter_pipeline_001:out_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [113:0] limiter_pipeline_001_source0_data;                                                                // limiter_pipeline_001:out_data -> limiter:rsp_sink_data
	wire   [24:0] limiter_pipeline_001_source0_channel;                                                             // limiter_pipeline_001:out_channel -> limiter:rsp_sink_channel
	wire          limiter_pipeline_001_source0_ready;                                                               // limiter:rsp_sink_ready -> limiter_pipeline_001:out_ready
	wire          cmd_xbar_demux_src0_ready;                                                                        // agent_pipeline:in_ready -> cmd_xbar_demux:src0_ready
	wire          agent_pipeline_source0_endofpacket;                                                               // agent_pipeline:out_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_source0_valid;                                                                     // agent_pipeline:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_source0_startofpacket;                                                             // agent_pipeline:out_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [113:0] agent_pipeline_source0_data;                                                                      // agent_pipeline:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [24:0] agent_pipeline_source0_channel;                                                                   // agent_pipeline:out_channel -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_source0_ready;                                                                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline:out_ready
	wire          agent_pipeline_001_source0_endofpacket;                                                           // agent_pipeline_001:out_endofpacket -> id_router:sink_endofpacket
	wire          agent_pipeline_001_source0_valid;                                                                 // agent_pipeline_001:out_valid -> id_router:sink_valid
	wire          agent_pipeline_001_source0_startofpacket;                                                         // agent_pipeline_001:out_startofpacket -> id_router:sink_startofpacket
	wire  [113:0] agent_pipeline_001_source0_data;                                                                  // agent_pipeline_001:out_data -> id_router:sink_data
	wire          agent_pipeline_001_source0_ready;                                                                 // id_router:sink_ready -> agent_pipeline_001:out_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_001:in_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_001:in_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_001:in_startofpacket
	wire  [113:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_001:in_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // agent_pipeline_001:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cmd_xbar_demux_src1_ready;                                                                        // agent_pipeline_002:in_ready -> cmd_xbar_demux:src1_ready
	wire          agent_pipeline_002_source0_endofpacket;                                                           // agent_pipeline_002:out_endofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_002_source0_valid;                                                                 // agent_pipeline_002:out_valid -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_002_source0_startofpacket;                                                         // agent_pipeline_002:out_startofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [113:0] agent_pipeline_002_source0_data;                                                                  // agent_pipeline_002:out_data -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [24:0] agent_pipeline_002_source0_channel;                                                               // agent_pipeline_002:out_channel -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_002_source0_ready;                                                                 // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_002:out_ready
	wire          agent_pipeline_003_source0_endofpacket;                                                           // agent_pipeline_003:out_endofpacket -> id_router_001:sink_endofpacket
	wire          agent_pipeline_003_source0_valid;                                                                 // agent_pipeline_003:out_valid -> id_router_001:sink_valid
	wire          agent_pipeline_003_source0_startofpacket;                                                         // agent_pipeline_003:out_startofpacket -> id_router_001:sink_startofpacket
	wire  [113:0] agent_pipeline_003_source0_data;                                                                  // agent_pipeline_003:out_data -> id_router_001:sink_data
	wire          agent_pipeline_003_source0_ready;                                                                 // id_router_001:sink_ready -> agent_pipeline_003:out_ready
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_003:in_endofpacket
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                      // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_003:in_valid
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;              // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_003:in_startofpacket
	wire  [113:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                       // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_003:in_data
	wire          sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                      // agent_pipeline_003:in_ready -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cmd_xbar_demux_src2_ready;                                                                        // agent_pipeline_004:in_ready -> cmd_xbar_demux:src2_ready
	wire          agent_pipeline_004_source0_endofpacket;                                                           // agent_pipeline_004:out_endofpacket -> audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_004_source0_valid;                                                                 // agent_pipeline_004:out_valid -> audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_004_source0_startofpacket;                                                         // agent_pipeline_004:out_startofpacket -> audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [113:0] agent_pipeline_004_source0_data;                                                                  // agent_pipeline_004:out_data -> audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [24:0] agent_pipeline_004_source0_channel;                                                               // agent_pipeline_004:out_channel -> audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_004_source0_ready;                                                                 // audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_004:out_ready
	wire          agent_pipeline_005_source0_endofpacket;                                                           // agent_pipeline_005:out_endofpacket -> id_router_002:sink_endofpacket
	wire          agent_pipeline_005_source0_valid;                                                                 // agent_pipeline_005:out_valid -> id_router_002:sink_valid
	wire          agent_pipeline_005_source0_startofpacket;                                                         // agent_pipeline_005:out_startofpacket -> id_router_002:sink_startofpacket
	wire  [113:0] agent_pipeline_005_source0_data;                                                                  // agent_pipeline_005:out_data -> id_router_002:sink_data
	wire          agent_pipeline_005_source0_ready;                                                                 // id_router_002:sink_ready -> agent_pipeline_005:out_ready
	wire          audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                    // audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_005:in_endofpacket
	wire          audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rp_valid;                          // audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_005:in_valid
	wire          audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                  // audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_005:in_startofpacket
	wire  [113:0] audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rp_data;                           // audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_005:in_data
	wire          audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rp_ready;                          // agent_pipeline_005:in_ready -> audio_data_fregen_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cmd_xbar_demux_src3_ready;                                                                        // agent_pipeline_006:in_ready -> cmd_xbar_demux:src3_ready
	wire          agent_pipeline_006_source0_endofpacket;                                                           // agent_pipeline_006:out_endofpacket -> audio_empty_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_006_source0_valid;                                                                 // agent_pipeline_006:out_valid -> audio_empty_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_006_source0_startofpacket;                                                         // agent_pipeline_006:out_startofpacket -> audio_empty_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [113:0] agent_pipeline_006_source0_data;                                                                  // agent_pipeline_006:out_data -> audio_empty_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [24:0] agent_pipeline_006_source0_channel;                                                               // agent_pipeline_006:out_channel -> audio_empty_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_006_source0_ready;                                                                 // audio_empty_s1_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_006:out_ready
	wire          agent_pipeline_007_source0_endofpacket;                                                           // agent_pipeline_007:out_endofpacket -> id_router_003:sink_endofpacket
	wire          agent_pipeline_007_source0_valid;                                                                 // agent_pipeline_007:out_valid -> id_router_003:sink_valid
	wire          agent_pipeline_007_source0_startofpacket;                                                         // agent_pipeline_007:out_startofpacket -> id_router_003:sink_startofpacket
	wire  [113:0] agent_pipeline_007_source0_data;                                                                  // agent_pipeline_007:out_data -> id_router_003:sink_data
	wire          agent_pipeline_007_source0_ready;                                                                 // id_router_003:sink_ready -> agent_pipeline_007:out_ready
	wire          audio_empty_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                          // audio_empty_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_007:in_endofpacket
	wire          audio_empty_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                // audio_empty_s1_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_007:in_valid
	wire          audio_empty_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                        // audio_empty_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_007:in_startofpacket
	wire  [113:0] audio_empty_s1_translator_avalon_universal_slave_0_agent_rp_data;                                 // audio_empty_s1_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_007:in_data
	wire          audio_empty_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                // agent_pipeline_007:in_ready -> audio_empty_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cmd_xbar_demux_src4_ready;                                                                        // agent_pipeline_008:in_ready -> cmd_xbar_demux:src4_ready
	wire          agent_pipeline_008_source0_endofpacket;                                                           // agent_pipeline_008:out_endofpacket -> audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_008_source0_valid;                                                                 // agent_pipeline_008:out_valid -> audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_008_source0_startofpacket;                                                         // agent_pipeline_008:out_startofpacket -> audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [113:0] agent_pipeline_008_source0_data;                                                                  // agent_pipeline_008:out_data -> audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [24:0] agent_pipeline_008_source0_channel;                                                               // agent_pipeline_008:out_channel -> audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_008_source0_ready;                                                                 // audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_008:out_ready
	wire          agent_pipeline_009_source0_endofpacket;                                                           // agent_pipeline_009:out_endofpacket -> id_router_004:sink_endofpacket
	wire          agent_pipeline_009_source0_valid;                                                                 // agent_pipeline_009:out_valid -> id_router_004:sink_valid
	wire          agent_pipeline_009_source0_startofpacket;                                                         // agent_pipeline_009:out_startofpacket -> id_router_004:sink_startofpacket
	wire  [113:0] agent_pipeline_009_source0_data;                                                                  // agent_pipeline_009:out_data -> id_router_004:sink_data
	wire          agent_pipeline_009_source0_ready;                                                                 // id_router_004:sink_ready -> agent_pipeline_009:out_ready
	wire          audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_009:in_endofpacket
	wire          audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rp_valid;                            // audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_009:in_valid
	wire          audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_009:in_startofpacket
	wire  [113:0] audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rp_data;                             // audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_009:in_data
	wire          audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rp_ready;                            // agent_pipeline_009:in_ready -> audio_fifo_full_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cmd_xbar_demux_src5_ready;                                                                        // agent_pipeline_010:in_ready -> cmd_xbar_demux:src5_ready
	wire          agent_pipeline_010_source0_endofpacket;                                                           // agent_pipeline_010:out_endofpacket -> audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_010_source0_valid;                                                                 // agent_pipeline_010:out_valid -> audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_010_source0_startofpacket;                                                         // agent_pipeline_010:out_startofpacket -> audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [113:0] agent_pipeline_010_source0_data;                                                                  // agent_pipeline_010:out_data -> audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [24:0] agent_pipeline_010_source0_channel;                                                               // agent_pipeline_010:out_channel -> audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_010_source0_ready;                                                                 // audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_010:out_ready
	wire          agent_pipeline_011_source0_endofpacket;                                                           // agent_pipeline_011:out_endofpacket -> id_router_005:sink_endofpacket
	wire          agent_pipeline_011_source0_valid;                                                                 // agent_pipeline_011:out_valid -> id_router_005:sink_valid
	wire          agent_pipeline_011_source0_startofpacket;                                                         // agent_pipeline_011:out_startofpacket -> id_router_005:sink_startofpacket
	wire  [113:0] agent_pipeline_011_source0_data;                                                                  // agent_pipeline_011:out_data -> id_router_005:sink_data
	wire          agent_pipeline_011_source0_ready;                                                                 // id_router_005:sink_ready -> agent_pipeline_011:out_ready
	wire          audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_011:in_endofpacket
	wire          audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rp_valid;                            // audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_011:in_valid
	wire          audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_011:in_startofpacket
	wire  [113:0] audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rp_data;                             // audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_011:in_data
	wire          audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rp_ready;                            // agent_pipeline_011:in_ready -> audio_fifo_used_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cmd_xbar_mux_006_src_endofpacket;                                                                 // cmd_xbar_mux_006:src_endofpacket -> agent_pipeline_012:in_endofpacket
	wire          cmd_xbar_mux_006_src_valid;                                                                       // cmd_xbar_mux_006:src_valid -> agent_pipeline_012:in_valid
	wire          cmd_xbar_mux_006_src_startofpacket;                                                               // cmd_xbar_mux_006:src_startofpacket -> agent_pipeline_012:in_startofpacket
	wire  [113:0] cmd_xbar_mux_006_src_data;                                                                        // cmd_xbar_mux_006:src_data -> agent_pipeline_012:in_data
	wire   [24:0] cmd_xbar_mux_006_src_channel;                                                                     // cmd_xbar_mux_006:src_channel -> agent_pipeline_012:in_channel
	wire          cmd_xbar_mux_006_src_ready;                                                                       // agent_pipeline_012:in_ready -> cmd_xbar_mux_006:src_ready
	wire          agent_pipeline_012_source0_endofpacket;                                                           // agent_pipeline_012:out_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_012_source0_valid;                                                                 // agent_pipeline_012:out_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_012_source0_startofpacket;                                                         // agent_pipeline_012:out_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [113:0] agent_pipeline_012_source0_data;                                                                  // agent_pipeline_012:out_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [24:0] agent_pipeline_012_source0_channel;                                                               // agent_pipeline_012:out_channel -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_012_source0_ready;                                                                 // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_012:out_ready
	wire          agent_pipeline_013_source0_endofpacket;                                                           // agent_pipeline_013:out_endofpacket -> id_router_006:sink_endofpacket
	wire          agent_pipeline_013_source0_valid;                                                                 // agent_pipeline_013:out_valid -> id_router_006:sink_valid
	wire          agent_pipeline_013_source0_startofpacket;                                                         // agent_pipeline_013:out_startofpacket -> id_router_006:sink_startofpacket
	wire  [113:0] agent_pipeline_013_source0_data;                                                                  // agent_pipeline_013:out_data -> id_router_006:sink_data
	wire          agent_pipeline_013_source0_ready;                                                                 // id_router_006:sink_ready -> agent_pipeline_013:out_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_013:in_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                         // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_013:in_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_013:in_startofpacket
	wire  [113:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                          // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_013:in_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                         // agent_pipeline_013:in_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cmd_xbar_demux_src7_ready;                                                                        // agent_pipeline_014:in_ready -> cmd_xbar_demux:src7_ready
	wire          agent_pipeline_014_source0_endofpacket;                                                           // agent_pipeline_014:out_endofpacket -> audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_014_source0_valid;                                                                 // agent_pipeline_014:out_valid -> audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_014_source0_startofpacket;                                                         // agent_pipeline_014:out_startofpacket -> audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [113:0] agent_pipeline_014_source0_data;                                                                  // agent_pipeline_014:out_data -> audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [24:0] agent_pipeline_014_source0_channel;                                                               // agent_pipeline_014:out_channel -> audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_014_source0_ready;                                                                 // audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_014:out_ready
	wire          agent_pipeline_015_source0_endofpacket;                                                           // agent_pipeline_015:out_endofpacket -> id_router_007:sink_endofpacket
	wire          agent_pipeline_015_source0_valid;                                                                 // agent_pipeline_015:out_valid -> id_router_007:sink_valid
	wire          agent_pipeline_015_source0_startofpacket;                                                         // agent_pipeline_015:out_startofpacket -> id_router_007:sink_startofpacket
	wire  [113:0] agent_pipeline_015_source0_data;                                                                  // agent_pipeline_015:out_data -> id_router_007:sink_data
	wire          agent_pipeline_015_source0_ready;                                                                 // id_router_007:sink_ready -> agent_pipeline_015:out_ready
	wire          audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                 // audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_015:in_endofpacket
	wire          audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rp_valid;                       // audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_015:in_valid
	wire          audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;               // audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_015:in_startofpacket
	wire  [113:0] audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rp_data;                        // audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_015:in_data
	wire          audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rp_ready;                       // agent_pipeline_015:in_ready -> audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cmd_xbar_demux_src8_ready;                                                                        // agent_pipeline_016:in_ready -> cmd_xbar_demux:src8_ready
	wire          agent_pipeline_016_source0_endofpacket;                                                           // agent_pipeline_016:out_endofpacket -> audio_out_pause_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_016_source0_valid;                                                                 // agent_pipeline_016:out_valid -> audio_out_pause_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_016_source0_startofpacket;                                                         // agent_pipeline_016:out_startofpacket -> audio_out_pause_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [113:0] agent_pipeline_016_source0_data;                                                                  // agent_pipeline_016:out_data -> audio_out_pause_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [24:0] agent_pipeline_016_source0_channel;                                                               // agent_pipeline_016:out_channel -> audio_out_pause_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_016_source0_ready;                                                                 // audio_out_pause_s1_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_016:out_ready
	wire          agent_pipeline_017_source0_endofpacket;                                                           // agent_pipeline_017:out_endofpacket -> id_router_008:sink_endofpacket
	wire          agent_pipeline_017_source0_valid;                                                                 // agent_pipeline_017:out_valid -> id_router_008:sink_valid
	wire          agent_pipeline_017_source0_startofpacket;                                                         // agent_pipeline_017:out_startofpacket -> id_router_008:sink_startofpacket
	wire  [113:0] agent_pipeline_017_source0_data;                                                                  // agent_pipeline_017:out_data -> id_router_008:sink_data
	wire          agent_pipeline_017_source0_ready;                                                                 // id_router_008:sink_ready -> agent_pipeline_017:out_ready
	wire          audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // audio_out_pause_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_017:in_endofpacket
	wire          audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rp_valid;                            // audio_out_pause_s1_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_017:in_valid
	wire          audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // audio_out_pause_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_017:in_startofpacket
	wire  [113:0] audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rp_data;                             // audio_out_pause_s1_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_017:in_data
	wire          audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rp_ready;                            // agent_pipeline_017:in_ready -> audio_out_pause_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cmd_xbar_demux_src9_ready;                                                                        // agent_pipeline_018:in_ready -> cmd_xbar_demux:src9_ready
	wire          agent_pipeline_018_source0_endofpacket;                                                           // agent_pipeline_018:out_endofpacket -> audio_out_stop_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_018_source0_valid;                                                                 // agent_pipeline_018:out_valid -> audio_out_stop_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_018_source0_startofpacket;                                                         // agent_pipeline_018:out_startofpacket -> audio_out_stop_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [113:0] agent_pipeline_018_source0_data;                                                                  // agent_pipeline_018:out_data -> audio_out_stop_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [24:0] agent_pipeline_018_source0_channel;                                                               // agent_pipeline_018:out_channel -> audio_out_stop_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_018_source0_ready;                                                                 // audio_out_stop_s1_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_018:out_ready
	wire          agent_pipeline_019_source0_endofpacket;                                                           // agent_pipeline_019:out_endofpacket -> id_router_009:sink_endofpacket
	wire          agent_pipeline_019_source0_valid;                                                                 // agent_pipeline_019:out_valid -> id_router_009:sink_valid
	wire          agent_pipeline_019_source0_startofpacket;                                                         // agent_pipeline_019:out_startofpacket -> id_router_009:sink_startofpacket
	wire  [113:0] agent_pipeline_019_source0_data;                                                                  // agent_pipeline_019:out_data -> id_router_009:sink_data
	wire          agent_pipeline_019_source0_ready;                                                                 // id_router_009:sink_ready -> agent_pipeline_019:out_ready
	wire          audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // audio_out_stop_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_019:in_endofpacket
	wire          audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rp_valid;                             // audio_out_stop_s1_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_019:in_valid
	wire          audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // audio_out_stop_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_019:in_startofpacket
	wire  [113:0] audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rp_data;                              // audio_out_stop_s1_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_019:in_data
	wire          audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rp_ready;                             // agent_pipeline_019:in_ready -> audio_out_stop_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cmd_xbar_demux_src10_ready;                                                                       // agent_pipeline_020:in_ready -> cmd_xbar_demux:src10_ready
	wire          agent_pipeline_020_source0_endofpacket;                                                           // agent_pipeline_020:out_endofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_020_source0_valid;                                                                 // agent_pipeline_020:out_valid -> timer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_020_source0_startofpacket;                                                         // agent_pipeline_020:out_startofpacket -> timer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [113:0] agent_pipeline_020_source0_data;                                                                  // agent_pipeline_020:out_data -> timer_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [24:0] agent_pipeline_020_source0_channel;                                                               // agent_pipeline_020:out_channel -> timer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_020_source0_ready;                                                                 // timer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_020:out_ready
	wire          agent_pipeline_021_source0_endofpacket;                                                           // agent_pipeline_021:out_endofpacket -> id_router_010:sink_endofpacket
	wire          agent_pipeline_021_source0_valid;                                                                 // agent_pipeline_021:out_valid -> id_router_010:sink_valid
	wire          agent_pipeline_021_source0_startofpacket;                                                         // agent_pipeline_021:out_startofpacket -> id_router_010:sink_startofpacket
	wire  [113:0] agent_pipeline_021_source0_data;                                                                  // agent_pipeline_021:out_data -> id_router_010:sink_data
	wire          agent_pipeline_021_source0_ready;                                                                 // id_router_010:sink_ready -> agent_pipeline_021:out_ready
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // timer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_021:in_endofpacket
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // timer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_021:in_valid
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // timer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_021:in_startofpacket
	wire  [113:0] timer_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // timer_s1_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_021:in_data
	wire          timer_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // agent_pipeline_021:in_ready -> timer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cmd_xbar_demux_src11_ready;                                                                       // agent_pipeline_022:in_ready -> cmd_xbar_demux:src11_ready
	wire          agent_pipeline_022_source0_endofpacket;                                                           // agent_pipeline_022:out_endofpacket -> key_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_022_source0_valid;                                                                 // agent_pipeline_022:out_valid -> key_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_022_source0_startofpacket;                                                         // agent_pipeline_022:out_startofpacket -> key_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [113:0] agent_pipeline_022_source0_data;                                                                  // agent_pipeline_022:out_data -> key_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [24:0] agent_pipeline_022_source0_channel;                                                               // agent_pipeline_022:out_channel -> key_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_022_source0_ready;                                                                 // key_s1_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_022:out_ready
	wire          agent_pipeline_023_source0_endofpacket;                                                           // agent_pipeline_023:out_endofpacket -> id_router_011:sink_endofpacket
	wire          agent_pipeline_023_source0_valid;                                                                 // agent_pipeline_023:out_valid -> id_router_011:sink_valid
	wire          agent_pipeline_023_source0_startofpacket;                                                         // agent_pipeline_023:out_startofpacket -> id_router_011:sink_startofpacket
	wire  [113:0] agent_pipeline_023_source0_data;                                                                  // agent_pipeline_023:out_data -> id_router_011:sink_data
	wire          agent_pipeline_023_source0_ready;                                                                 // id_router_011:sink_ready -> agent_pipeline_023:out_ready
	wire          key_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // key_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_023:in_endofpacket
	wire          key_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // key_s1_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_023:in_valid
	wire          key_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // key_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_023:in_startofpacket
	wire  [113:0] key_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // key_s1_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_023:in_data
	wire          key_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // agent_pipeline_023:in_ready -> key_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cmd_xbar_demux_src12_ready;                                                                       // agent_pipeline_024:in_ready -> cmd_xbar_demux:src12_ready
	wire          agent_pipeline_024_source0_endofpacket;                                                           // agent_pipeline_024:out_endofpacket -> signal_selector_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_024_source0_valid;                                                                 // agent_pipeline_024:out_valid -> signal_selector_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_024_source0_startofpacket;                                                         // agent_pipeline_024:out_startofpacket -> signal_selector_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [113:0] agent_pipeline_024_source0_data;                                                                  // agent_pipeline_024:out_data -> signal_selector_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [24:0] agent_pipeline_024_source0_channel;                                                               // agent_pipeline_024:out_channel -> signal_selector_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_024_source0_ready;                                                                 // signal_selector_s1_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_024:out_ready
	wire          agent_pipeline_025_source0_endofpacket;                                                           // agent_pipeline_025:out_endofpacket -> id_router_012:sink_endofpacket
	wire          agent_pipeline_025_source0_valid;                                                                 // agent_pipeline_025:out_valid -> id_router_012:sink_valid
	wire          agent_pipeline_025_source0_startofpacket;                                                         // agent_pipeline_025:out_startofpacket -> id_router_012:sink_startofpacket
	wire  [113:0] agent_pipeline_025_source0_data;                                                                  // agent_pipeline_025:out_data -> id_router_012:sink_data
	wire          agent_pipeline_025_source0_ready;                                                                 // id_router_012:sink_ready -> agent_pipeline_025:out_ready
	wire          signal_selector_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // signal_selector_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_025:in_endofpacket
	wire          signal_selector_s1_translator_avalon_universal_slave_0_agent_rp_valid;                            // signal_selector_s1_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_025:in_valid
	wire          signal_selector_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // signal_selector_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_025:in_startofpacket
	wire  [113:0] signal_selector_s1_translator_avalon_universal_slave_0_agent_rp_data;                             // signal_selector_s1_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_025:in_data
	wire          signal_selector_s1_translator_avalon_universal_slave_0_agent_rp_ready;                            // agent_pipeline_025:in_ready -> signal_selector_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cmd_xbar_demux_src13_ready;                                                                       // agent_pipeline_026:in_ready -> cmd_xbar_demux:src13_ready
	wire          agent_pipeline_026_source0_endofpacket;                                                           // agent_pipeline_026:out_endofpacket -> modulation_selector_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_026_source0_valid;                                                                 // agent_pipeline_026:out_valid -> modulation_selector_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_026_source0_startofpacket;                                                         // agent_pipeline_026:out_startofpacket -> modulation_selector_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [113:0] agent_pipeline_026_source0_data;                                                                  // agent_pipeline_026:out_data -> modulation_selector_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [24:0] agent_pipeline_026_source0_channel;                                                               // agent_pipeline_026:out_channel -> modulation_selector_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_026_source0_ready;                                                                 // modulation_selector_s1_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_026:out_ready
	wire          agent_pipeline_027_source0_endofpacket;                                                           // agent_pipeline_027:out_endofpacket -> id_router_013:sink_endofpacket
	wire          agent_pipeline_027_source0_valid;                                                                 // agent_pipeline_027:out_valid -> id_router_013:sink_valid
	wire          agent_pipeline_027_source0_startofpacket;                                                         // agent_pipeline_027:out_startofpacket -> id_router_013:sink_startofpacket
	wire  [113:0] agent_pipeline_027_source0_data;                                                                  // agent_pipeline_027:out_data -> id_router_013:sink_data
	wire          agent_pipeline_027_source0_ready;                                                                 // id_router_013:sink_ready -> agent_pipeline_027:out_ready
	wire          modulation_selector_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                  // modulation_selector_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_027:in_endofpacket
	wire          modulation_selector_s1_translator_avalon_universal_slave_0_agent_rp_valid;                        // modulation_selector_s1_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_027:in_valid
	wire          modulation_selector_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                // modulation_selector_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_027:in_startofpacket
	wire  [113:0] modulation_selector_s1_translator_avalon_universal_slave_0_agent_rp_data;                         // modulation_selector_s1_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_027:in_data
	wire          modulation_selector_s1_translator_avalon_universal_slave_0_agent_rp_ready;                        // agent_pipeline_027:in_ready -> modulation_selector_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          crosser_out_ready;                                                                                // agent_pipeline_028:in_ready -> crosser:out_ready
	wire          agent_pipeline_028_source0_endofpacket;                                                           // agent_pipeline_028:out_endofpacket -> keyboard_keys_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_028_source0_valid;                                                                 // agent_pipeline_028:out_valid -> keyboard_keys_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_028_source0_startofpacket;                                                         // agent_pipeline_028:out_startofpacket -> keyboard_keys_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [113:0] agent_pipeline_028_source0_data;                                                                  // agent_pipeline_028:out_data -> keyboard_keys_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [24:0] agent_pipeline_028_source0_channel;                                                               // agent_pipeline_028:out_channel -> keyboard_keys_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_028_source0_ready;                                                                 // keyboard_keys_s1_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_028:out_ready
	wire          agent_pipeline_029_source0_endofpacket;                                                           // agent_pipeline_029:out_endofpacket -> id_router_014:sink_endofpacket
	wire          agent_pipeline_029_source0_valid;                                                                 // agent_pipeline_029:out_valid -> id_router_014:sink_valid
	wire          agent_pipeline_029_source0_startofpacket;                                                         // agent_pipeline_029:out_startofpacket -> id_router_014:sink_startofpacket
	wire  [113:0] agent_pipeline_029_source0_data;                                                                  // agent_pipeline_029:out_data -> id_router_014:sink_data
	wire          agent_pipeline_029_source0_ready;                                                                 // id_router_014:sink_ready -> agent_pipeline_029:out_ready
	wire          keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // keyboard_keys_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_029:in_endofpacket
	wire          keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rp_valid;                              // keyboard_keys_s1_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_029:in_valid
	wire          keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // keyboard_keys_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_029:in_startofpacket
	wire  [113:0] keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rp_data;                               // keyboard_keys_s1_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_029:in_data
	wire          keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rp_ready;                              // agent_pipeline_029:in_ready -> keyboard_keys_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          crosser_001_out_ready;                                                                            // agent_pipeline_030:in_ready -> crosser_001:out_ready
	wire          agent_pipeline_030_source0_endofpacket;                                                           // agent_pipeline_030:out_endofpacket -> mouse_pos_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_030_source0_valid;                                                                 // agent_pipeline_030:out_valid -> mouse_pos_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_030_source0_startofpacket;                                                         // agent_pipeline_030:out_startofpacket -> mouse_pos_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [113:0] agent_pipeline_030_source0_data;                                                                  // agent_pipeline_030:out_data -> mouse_pos_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [24:0] agent_pipeline_030_source0_channel;                                                               // agent_pipeline_030:out_channel -> mouse_pos_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_030_source0_ready;                                                                 // mouse_pos_s1_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_030:out_ready
	wire          agent_pipeline_031_source0_endofpacket;                                                           // agent_pipeline_031:out_endofpacket -> id_router_015:sink_endofpacket
	wire          agent_pipeline_031_source0_valid;                                                                 // agent_pipeline_031:out_valid -> id_router_015:sink_valid
	wire          agent_pipeline_031_source0_startofpacket;                                                         // agent_pipeline_031:out_startofpacket -> id_router_015:sink_startofpacket
	wire  [113:0] agent_pipeline_031_source0_data;                                                                  // agent_pipeline_031:out_data -> id_router_015:sink_data
	wire          agent_pipeline_031_source0_ready;                                                                 // id_router_015:sink_ready -> agent_pipeline_031:out_ready
	wire          mouse_pos_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // mouse_pos_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_031:in_endofpacket
	wire          mouse_pos_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // mouse_pos_s1_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_031:in_valid
	wire          mouse_pos_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // mouse_pos_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_031:in_startofpacket
	wire  [113:0] mouse_pos_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // mouse_pos_s1_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_031:in_data
	wire          mouse_pos_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // agent_pipeline_031:in_ready -> mouse_pos_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cmd_xbar_demux_src16_ready;                                                                       // agent_pipeline_032:in_ready -> cmd_xbar_demux:src16_ready
	wire          agent_pipeline_032_source0_endofpacket;                                                           // agent_pipeline_032:out_endofpacket -> div_freq_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_032_source0_valid;                                                                 // agent_pipeline_032:out_valid -> div_freq_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_032_source0_startofpacket;                                                         // agent_pipeline_032:out_startofpacket -> div_freq_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [113:0] agent_pipeline_032_source0_data;                                                                  // agent_pipeline_032:out_data -> div_freq_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [24:0] agent_pipeline_032_source0_channel;                                                               // agent_pipeline_032:out_channel -> div_freq_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_032_source0_ready;                                                                 // div_freq_s1_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_032:out_ready
	wire          agent_pipeline_033_source0_endofpacket;                                                           // agent_pipeline_033:out_endofpacket -> id_router_016:sink_endofpacket
	wire          agent_pipeline_033_source0_valid;                                                                 // agent_pipeline_033:out_valid -> id_router_016:sink_valid
	wire          agent_pipeline_033_source0_startofpacket;                                                         // agent_pipeline_033:out_startofpacket -> id_router_016:sink_startofpacket
	wire  [113:0] agent_pipeline_033_source0_data;                                                                  // agent_pipeline_033:out_data -> id_router_016:sink_data
	wire          agent_pipeline_033_source0_ready;                                                                 // id_router_016:sink_ready -> agent_pipeline_033:out_ready
	wire          div_freq_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // div_freq_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_033:in_endofpacket
	wire          div_freq_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                   // div_freq_s1_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_033:in_valid
	wire          div_freq_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // div_freq_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_033:in_startofpacket
	wire  [113:0] div_freq_s1_translator_avalon_universal_slave_0_agent_rp_data;                                    // div_freq_s1_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_033:in_data
	wire          div_freq_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                   // agent_pipeline_033:in_ready -> div_freq_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cmd_xbar_demux_src17_ready;                                                                       // agent_pipeline_034:in_ready -> cmd_xbar_demux:src17_ready
	wire          agent_pipeline_034_source0_endofpacket;                                                           // agent_pipeline_034:out_endofpacket -> audio_sel_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_034_source0_valid;                                                                 // agent_pipeline_034:out_valid -> audio_sel_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_034_source0_startofpacket;                                                         // agent_pipeline_034:out_startofpacket -> audio_sel_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [113:0] agent_pipeline_034_source0_data;                                                                  // agent_pipeline_034:out_data -> audio_sel_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [24:0] agent_pipeline_034_source0_channel;                                                               // agent_pipeline_034:out_channel -> audio_sel_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_034_source0_ready;                                                                 // audio_sel_s1_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_034:out_ready
	wire          agent_pipeline_035_source0_endofpacket;                                                           // agent_pipeline_035:out_endofpacket -> id_router_017:sink_endofpacket
	wire          agent_pipeline_035_source0_valid;                                                                 // agent_pipeline_035:out_valid -> id_router_017:sink_valid
	wire          agent_pipeline_035_source0_startofpacket;                                                         // agent_pipeline_035:out_startofpacket -> id_router_017:sink_startofpacket
	wire  [113:0] agent_pipeline_035_source0_data;                                                                  // agent_pipeline_035:out_data -> id_router_017:sink_data
	wire          agent_pipeline_035_source0_ready;                                                                 // id_router_017:sink_ready -> agent_pipeline_035:out_ready
	wire          audio_sel_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // audio_sel_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_035:in_endofpacket
	wire          audio_sel_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // audio_sel_s1_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_035:in_valid
	wire          audio_sel_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // audio_sel_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_035:in_startofpacket
	wire  [113:0] audio_sel_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // audio_sel_s1_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_035:in_data
	wire          audio_sel_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // agent_pipeline_035:in_ready -> audio_sel_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          crosser_002_out_ready;                                                                            // agent_pipeline_036:in_ready -> crosser_002:out_ready
	wire          agent_pipeline_036_source0_endofpacket;                                                           // agent_pipeline_036:out_endofpacket -> vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_036_source0_valid;                                                                 // agent_pipeline_036:out_valid -> vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_036_source0_startofpacket;                                                         // agent_pipeline_036:out_startofpacket -> vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [113:0] agent_pipeline_036_source0_data;                                                                  // agent_pipeline_036:out_data -> vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:cp_data
	wire   [24:0] agent_pipeline_036_source0_channel;                                                               // agent_pipeline_036:out_channel -> vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_036_source0_ready;                                                                 // vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_036:out_ready
	wire          agent_pipeline_037_source0_endofpacket;                                                           // agent_pipeline_037:out_endofpacket -> id_router_018:sink_endofpacket
	wire          agent_pipeline_037_source0_valid;                                                                 // agent_pipeline_037:out_valid -> id_router_018:sink_valid
	wire          agent_pipeline_037_source0_startofpacket;                                                         // agent_pipeline_037:out_startofpacket -> id_router_018:sink_startofpacket
	wire  [113:0] agent_pipeline_037_source0_data;                                                                  // agent_pipeline_037:out_data -> id_router_018:sink_data
	wire          agent_pipeline_037_source0_ready;                                                                 // id_router_018:sink_ready -> agent_pipeline_037:out_ready
	wire          vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rp_endofpacket;                // vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_037:in_endofpacket
	wire          vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rp_valid;                      // vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_037:in_valid
	wire          vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rp_startofpacket;              // vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_037:in_startofpacket
	wire  [113:0] vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rp_data;                       // vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_037:in_data
	wire          vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rp_ready;                      // agent_pipeline_037:in_ready -> vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cmd_xbar_demux_src19_ready;                                                                       // agent_pipeline_038:in_ready -> cmd_xbar_demux:src19_ready
	wire          agent_pipeline_038_source0_endofpacket;                                                           // agent_pipeline_038:out_endofpacket -> audio_wrclk_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_038_source0_valid;                                                                 // agent_pipeline_038:out_valid -> audio_wrclk_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_038_source0_startofpacket;                                                         // agent_pipeline_038:out_startofpacket -> audio_wrclk_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [113:0] agent_pipeline_038_source0_data;                                                                  // agent_pipeline_038:out_data -> audio_wrclk_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [24:0] agent_pipeline_038_source0_channel;                                                               // agent_pipeline_038:out_channel -> audio_wrclk_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_038_source0_ready;                                                                 // audio_wrclk_s1_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_038:out_ready
	wire          agent_pipeline_039_source0_endofpacket;                                                           // agent_pipeline_039:out_endofpacket -> id_router_019:sink_endofpacket
	wire          agent_pipeline_039_source0_valid;                                                                 // agent_pipeline_039:out_valid -> id_router_019:sink_valid
	wire          agent_pipeline_039_source0_startofpacket;                                                         // agent_pipeline_039:out_startofpacket -> id_router_019:sink_startofpacket
	wire  [113:0] agent_pipeline_039_source0_data;                                                                  // agent_pipeline_039:out_data -> id_router_019:sink_data
	wire          agent_pipeline_039_source0_ready;                                                                 // id_router_019:sink_ready -> agent_pipeline_039:out_ready
	wire          audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                          // audio_wrclk_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_039:in_endofpacket
	wire          audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                // audio_wrclk_s1_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_039:in_valid
	wire          audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                        // audio_wrclk_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_039:in_startofpacket
	wire  [113:0] audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rp_data;                                 // audio_wrclk_s1_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_039:in_data
	wire          audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                // agent_pipeline_039:in_ready -> audio_wrclk_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cmd_xbar_demux_src20_ready;                                                                       // agent_pipeline_040:in_ready -> cmd_xbar_demux:src20_ready
	wire          agent_pipeline_040_source0_endofpacket;                                                           // agent_pipeline_040:out_endofpacket -> audio_wrreq_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_040_source0_valid;                                                                 // agent_pipeline_040:out_valid -> audio_wrreq_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_040_source0_startofpacket;                                                         // agent_pipeline_040:out_startofpacket -> audio_wrreq_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [113:0] agent_pipeline_040_source0_data;                                                                  // agent_pipeline_040:out_data -> audio_wrreq_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [24:0] agent_pipeline_040_source0_channel;                                                               // agent_pipeline_040:out_channel -> audio_wrreq_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_040_source0_ready;                                                                 // audio_wrreq_s1_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_040:out_ready
	wire          agent_pipeline_041_source0_endofpacket;                                                           // agent_pipeline_041:out_endofpacket -> id_router_020:sink_endofpacket
	wire          agent_pipeline_041_source0_valid;                                                                 // agent_pipeline_041:out_valid -> id_router_020:sink_valid
	wire          agent_pipeline_041_source0_startofpacket;                                                         // agent_pipeline_041:out_startofpacket -> id_router_020:sink_startofpacket
	wire  [113:0] agent_pipeline_041_source0_data;                                                                  // agent_pipeline_041:out_data -> id_router_020:sink_data
	wire          agent_pipeline_041_source0_ready;                                                                 // id_router_020:sink_ready -> agent_pipeline_041:out_ready
	wire          audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                          // audio_wrreq_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_041:in_endofpacket
	wire          audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                // audio_wrreq_s1_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_041:in_valid
	wire          audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                        // audio_wrreq_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_041:in_startofpacket
	wire  [113:0] audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rp_data;                                 // audio_wrreq_s1_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_041:in_data
	wire          audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                // agent_pipeline_041:in_ready -> audio_wrreq_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          burst_adapter_source0_endofpacket;                                                                // burst_adapter:source0_endofpacket -> agent_pipeline_042:in_endofpacket
	wire          burst_adapter_source0_valid;                                                                      // burst_adapter:source0_valid -> agent_pipeline_042:in_valid
	wire          burst_adapter_source0_startofpacket;                                                              // burst_adapter:source0_startofpacket -> agent_pipeline_042:in_startofpacket
	wire   [95:0] burst_adapter_source0_data;                                                                       // burst_adapter:source0_data -> agent_pipeline_042:in_data
	wire          burst_adapter_source0_ready;                                                                      // agent_pipeline_042:in_ready -> burst_adapter:source0_ready
	wire   [24:0] burst_adapter_source0_channel;                                                                    // burst_adapter:source0_channel -> agent_pipeline_042:in_channel
	wire          agent_pipeline_042_source0_endofpacket;                                                           // agent_pipeline_042:out_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_042_source0_valid;                                                                 // agent_pipeline_042:out_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_042_source0_startofpacket;                                                         // agent_pipeline_042:out_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [95:0] agent_pipeline_042_source0_data;                                                                  // agent_pipeline_042:out_data -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [24:0] agent_pipeline_042_source0_channel;                                                               // agent_pipeline_042:out_channel -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_042_source0_ready;                                                                 // sdram_s1_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_042:out_ready
	wire          agent_pipeline_043_source0_endofpacket;                                                           // agent_pipeline_043:out_endofpacket -> id_router_021:sink_endofpacket
	wire          agent_pipeline_043_source0_valid;                                                                 // agent_pipeline_043:out_valid -> id_router_021:sink_valid
	wire          agent_pipeline_043_source0_startofpacket;                                                         // agent_pipeline_043:out_startofpacket -> id_router_021:sink_startofpacket
	wire   [95:0] agent_pipeline_043_source0_data;                                                                  // agent_pipeline_043:out_data -> id_router_021:sink_data
	wire          agent_pipeline_043_source0_ready;                                                                 // id_router_021:sink_ready -> agent_pipeline_043:out_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // sdram_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_043:in_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // sdram_s1_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_043:in_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // sdram_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_043:in_startofpacket
	wire   [95:0] sdram_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // sdram_s1_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_043:in_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // agent_pipeline_043:in_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cmd_xbar_demux_src22_ready;                                                                       // agent_pipeline_044:in_ready -> cmd_xbar_demux:src22_ready
	wire          agent_pipeline_044_source0_endofpacket;                                                           // agent_pipeline_044:out_endofpacket -> lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_044_source0_valid;                                                                 // agent_pipeline_044:out_valid -> lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_044_source0_startofpacket;                                                         // agent_pipeline_044:out_startofpacket -> lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [113:0] agent_pipeline_044_source0_data;                                                                  // agent_pipeline_044:out_data -> lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [24:0] agent_pipeline_044_source0_channel;                                                               // agent_pipeline_044:out_channel -> lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_044_source0_ready;                                                                 // lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_044:out_ready
	wire          agent_pipeline_045_source0_endofpacket;                                                           // agent_pipeline_045:out_endofpacket -> id_router_022:sink_endofpacket
	wire          agent_pipeline_045_source0_valid;                                                                 // agent_pipeline_045:out_valid -> id_router_022:sink_valid
	wire          agent_pipeline_045_source0_startofpacket;                                                         // agent_pipeline_045:out_startofpacket -> id_router_022:sink_startofpacket
	wire  [113:0] agent_pipeline_045_source0_data;                                                                  // agent_pipeline_045:out_data -> id_router_022:sink_data
	wire          agent_pipeline_045_source0_ready;                                                                 // id_router_022:sink_ready -> agent_pipeline_045:out_ready
	wire          lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;               // lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_045:in_endofpacket
	wire          lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rp_valid;                     // lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_045:in_valid
	wire          lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;             // lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_045:in_startofpacket
	wire  [113:0] lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rp_data;                      // lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_045:in_data
	wire          lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rp_ready;                     // agent_pipeline_045:in_ready -> lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cmd_xbar_demux_src23_ready;                                                                       // agent_pipeline_046:in_ready -> cmd_xbar_demux:src23_ready
	wire          agent_pipeline_046_source0_endofpacket;                                                           // agent_pipeline_046:out_endofpacket -> lfsr_val_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_046_source0_valid;                                                                 // agent_pipeline_046:out_valid -> lfsr_val_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_046_source0_startofpacket;                                                         // agent_pipeline_046:out_startofpacket -> lfsr_val_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [113:0] agent_pipeline_046_source0_data;                                                                  // agent_pipeline_046:out_data -> lfsr_val_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [24:0] agent_pipeline_046_source0_channel;                                                               // agent_pipeline_046:out_channel -> lfsr_val_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_046_source0_ready;                                                                 // lfsr_val_s1_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_046:out_ready
	wire          agent_pipeline_047_source0_endofpacket;                                                           // agent_pipeline_047:out_endofpacket -> id_router_023:sink_endofpacket
	wire          agent_pipeline_047_source0_valid;                                                                 // agent_pipeline_047:out_valid -> id_router_023:sink_valid
	wire          agent_pipeline_047_source0_startofpacket;                                                         // agent_pipeline_047:out_startofpacket -> id_router_023:sink_startofpacket
	wire  [113:0] agent_pipeline_047_source0_data;                                                                  // agent_pipeline_047:out_data -> id_router_023:sink_data
	wire          agent_pipeline_047_source0_ready;                                                                 // id_router_023:sink_ready -> agent_pipeline_047:out_ready
	wire          lfsr_val_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // lfsr_val_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_047:in_endofpacket
	wire          lfsr_val_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                   // lfsr_val_s1_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_047:in_valid
	wire          lfsr_val_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // lfsr_val_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_047:in_startofpacket
	wire  [113:0] lfsr_val_s1_translator_avalon_universal_slave_0_agent_rp_data;                                    // lfsr_val_s1_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_047:in_data
	wire          lfsr_val_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                   // agent_pipeline_047:in_ready -> lfsr_val_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cmd_xbar_demux_src24_ready;                                                                       // agent_pipeline_048:in_ready -> cmd_xbar_demux:src24_ready
	wire          agent_pipeline_048_source0_endofpacket;                                                           // agent_pipeline_048:out_endofpacket -> dds_increment_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          agent_pipeline_048_source0_valid;                                                                 // agent_pipeline_048:out_valid -> dds_increment_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          agent_pipeline_048_source0_startofpacket;                                                         // agent_pipeline_048:out_startofpacket -> dds_increment_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [113:0] agent_pipeline_048_source0_data;                                                                  // agent_pipeline_048:out_data -> dds_increment_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [24:0] agent_pipeline_048_source0_channel;                                                               // agent_pipeline_048:out_channel -> dds_increment_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          agent_pipeline_048_source0_ready;                                                                 // dds_increment_s1_translator_avalon_universal_slave_0_agent:cp_ready -> agent_pipeline_048:out_ready
	wire          agent_pipeline_049_source0_endofpacket;                                                           // agent_pipeline_049:out_endofpacket -> id_router_024:sink_endofpacket
	wire          agent_pipeline_049_source0_valid;                                                                 // agent_pipeline_049:out_valid -> id_router_024:sink_valid
	wire          agent_pipeline_049_source0_startofpacket;                                                         // agent_pipeline_049:out_startofpacket -> id_router_024:sink_startofpacket
	wire  [113:0] agent_pipeline_049_source0_data;                                                                  // agent_pipeline_049:out_data -> id_router_024:sink_data
	wire          agent_pipeline_049_source0_ready;                                                                 // id_router_024:sink_ready -> agent_pipeline_049:out_ready
	wire          dds_increment_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // dds_increment_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> agent_pipeline_049:in_endofpacket
	wire          dds_increment_s1_translator_avalon_universal_slave_0_agent_rp_valid;                              // dds_increment_s1_translator_avalon_universal_slave_0_agent:rp_valid -> agent_pipeline_049:in_valid
	wire          dds_increment_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // dds_increment_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> agent_pipeline_049:in_startofpacket
	wire  [113:0] dds_increment_s1_translator_avalon_universal_slave_0_agent_rp_data;                               // dds_increment_s1_translator_avalon_universal_slave_0_agent:rp_data -> agent_pipeline_049:in_data
	wire          dds_increment_s1_translator_avalon_universal_slave_0_agent_rp_ready;                              // agent_pipeline_049:in_ready -> dds_increment_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          irq_mapper_receiver1_irq;                                                                         // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire          irq_mapper_receiver2_irq;                                                                         // timer:irq -> irq_mapper:receiver2_irq
	wire          irq_mapper_receiver3_irq;                                                                         // key:irq -> irq_mapper:receiver3_irq
	wire   [31:0] cpu_d_irq_irq;                                                                                    // irq_mapper:sender_irq -> cpu:d_irq
	wire          irq_mapper_receiver0_irq;                                                                         // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire    [0:0] irq_synchronizer_receiver_irq;                                                                    // vga:alt_vip_vfr_0_interrupt_sender_irq -> irq_synchronizer:receiver_irq

	DE2_QSYS_audio audio (
		.clk_clk                      (clk_clk),                                                           //               clk.clk
		.data_divfrec_export          (audio2fifo_0_data_divfrec_export),                                  //      data_divfrec.export
		.data_fregen_s1_address       (audio_data_fregen_s1_translator_avalon_anti_slave_0_address),       //    data_fregen_s1.address
		.data_fregen_s1_write_n       (~audio_data_fregen_s1_translator_avalon_anti_slave_0_write),        //                  .write_n
		.data_fregen_s1_writedata     (audio_data_fregen_s1_translator_avalon_anti_slave_0_writedata),     //                  .writedata
		.data_fregen_s1_chipselect    (audio_data_fregen_s1_translator_avalon_anti_slave_0_chipselect),    //                  .chipselect
		.data_fregen_s1_readdata      (audio_data_fregen_s1_translator_avalon_anti_slave_0_readdata),      //                  .readdata
		.empty_export                 (audio2fifo_0_empty_export),                                         //             empty.export
		.empty_s1_address             (audio_empty_s1_translator_avalon_anti_slave_0_address),             //          empty_s1.address
		.empty_s1_readdata            (audio_empty_s1_translator_avalon_anti_slave_0_readdata),            //                  .readdata
		.fifo_full_export             (audio2fifo_0_fifo_full_export),                                     //         fifo_full.export
		.fifo_full_s1_address         (audio_fifo_full_s1_translator_avalon_anti_slave_0_address),         //      fifo_full_s1.address
		.fifo_full_s1_readdata        (audio_fifo_full_s1_translator_avalon_anti_slave_0_readdata),        //                  .readdata
		.fifo_used_export             (audio2fifo_0_fifo_used_export),                                     //         fifo_used.export
		.fifo_used_s1_address         (audio_fifo_used_s1_translator_avalon_anti_slave_0_address),         //      fifo_used_s1.address
		.fifo_used_s1_readdata        (audio_fifo_used_s1_translator_avalon_anti_slave_0_readdata),        //                  .readdata
		.out_data_audio_export        (audio2fifo_0_out_data_audio_export),                                //    out_data_audio.export
		.out_data_audio_s1_address    (audio_out_data_audio_s1_translator_avalon_anti_slave_0_address),    // out_data_audio_s1.address
		.out_data_audio_s1_write_n    (~audio_out_data_audio_s1_translator_avalon_anti_slave_0_write),     //                  .write_n
		.out_data_audio_s1_writedata  (audio_out_data_audio_s1_translator_avalon_anti_slave_0_writedata),  //                  .writedata
		.out_data_audio_s1_chipselect (audio_out_data_audio_s1_translator_avalon_anti_slave_0_chipselect), //                  .chipselect
		.out_data_audio_s1_readdata   (audio_out_data_audio_s1_translator_avalon_anti_slave_0_readdata),   //                  .readdata
		.out_pause_export             (audio2fifo_0_out_pause_export),                                     //         out_pause.export
		.out_pause_s1_address         (audio_out_pause_s1_translator_avalon_anti_slave_0_address),         //      out_pause_s1.address
		.out_pause_s1_write_n         (~audio_out_pause_s1_translator_avalon_anti_slave_0_write),          //                  .write_n
		.out_pause_s1_writedata       (audio_out_pause_s1_translator_avalon_anti_slave_0_writedata),       //                  .writedata
		.out_pause_s1_chipselect      (audio_out_pause_s1_translator_avalon_anti_slave_0_chipselect),      //                  .chipselect
		.out_pause_s1_readdata        (audio_out_pause_s1_translator_avalon_anti_slave_0_readdata),        //                  .readdata
		.out_stop_export              (audio2fifo_0_out_stop_export),                                      //          out_stop.export
		.out_stop_s1_address          (audio_out_stop_s1_translator_avalon_anti_slave_0_address),          //       out_stop_s1.address
		.out_stop_s1_write_n          (~audio_out_stop_s1_translator_avalon_anti_slave_0_write),           //                  .write_n
		.out_stop_s1_writedata        (audio_out_stop_s1_translator_avalon_anti_slave_0_writedata),        //                  .writedata
		.out_stop_s1_chipselect       (audio_out_stop_s1_translator_avalon_anti_slave_0_chipselect),       //                  .chipselect
		.out_stop_s1_readdata         (audio_out_stop_s1_translator_avalon_anti_slave_0_readdata),         //                  .readdata
		.reset_reset_n                (~rst_controller_reset_out_reset),                                   //             reset.reset_n
		.wrclk_export                 (audio2fifo_0_wrclk_export),                                         //             wrclk.export
		.wrclk_s1_address             (audio_wrclk_s1_translator_avalon_anti_slave_0_address),             //          wrclk_s1.address
		.wrclk_s1_write_n             (~audio_wrclk_s1_translator_avalon_anti_slave_0_write),              //                  .write_n
		.wrclk_s1_writedata           (audio_wrclk_s1_translator_avalon_anti_slave_0_writedata),           //                  .writedata
		.wrclk_s1_chipselect          (audio_wrclk_s1_translator_avalon_anti_slave_0_chipselect),          //                  .chipselect
		.wrclk_s1_readdata            (audio_wrclk_s1_translator_avalon_anti_slave_0_readdata),            //                  .readdata
		.wrreq_export                 (audio2fifo_0_wrreq_export),                                         //             wrreq.export
		.wrreq_s1_address             (audio_wrreq_s1_translator_avalon_anti_slave_0_address),             //          wrreq_s1.address
		.wrreq_s1_write_n             (~audio_wrreq_s1_translator_avalon_anti_slave_0_write),              //                  .write_n
		.wrreq_s1_writedata           (audio_wrreq_s1_translator_avalon_anti_slave_0_writedata),           //                  .writedata
		.wrreq_s1_chipselect          (audio_wrreq_s1_translator_avalon_anti_slave_0_chipselect),          //                  .chipselect
		.wrreq_s1_readdata            (audio_wrreq_s1_translator_avalon_anti_slave_0_readdata)             //                  .readdata
	);

	DE2_QSYS_audio_sel audio_sel (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                        //               reset.reset_n
		.address    (audio_sel_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~audio_sel_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (audio_sel_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (audio_sel_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (audio_sel_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (audio_sel_export)                                        // external_connection.export
	);

	DE2_QSYS_cpu cpu (
		.clk                                   (clk_clk),                                                          //                       clk.clk
		.reset_n                               (~rst_controller_001_reset_out_reset),                              //                   reset_n.reset_n
		.d_address                             (cpu_data_master_address),                                          //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                                       //                          .byteenable
		.d_read                                (cpu_data_master_read),                                             //                          .read
		.d_readdata                            (cpu_data_master_readdata),                                         //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                                      //                          .waitrequest
		.d_write                               (cpu_data_master_write),                                            //                          .write
		.d_writedata                           (cpu_data_master_writedata),                                        //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                                      //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                                   //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                                      //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                                  //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                               //                          .waitrequest
		.i_readdatavalid                       (cpu_instruction_master_readdatavalid),                             //                          .readdatavalid
		.d_irq                                 (cpu_d_irq_irq),                                                    //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                                //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (cpu_jtag_debug_module_translator_avalon_anti_slave_0_read),        //                          .read
		.jtag_debug_module_readdata            (cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),       //                          .write
		.jtag_debug_module_writedata           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                                  // custom_instruction_master.readra
	);

	DE2_QSYS_div_freq div_freq (
		.clk        (clk_clk),                                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                       //               reset.reset_n
		.address    (div_freq_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~div_freq_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (div_freq_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (div_freq_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (div_freq_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (div_freq_export)                                        // external_connection.export
	);

	DE2_QSYS_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                                //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                        //             reset.reset_n
		.av_chipselect  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                                //               irq.irq
	);

	DE2_QSYS_key key (
		.clk        (clk_clk),                                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (key_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~key_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (key_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (key_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (key_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (key_external_connection_export),                   // external_connection.export
		.irq        (irq_mapper_receiver3_irq)                          //                 irq.irq
	);

	DE2_QSYS_keyboard_keys keyboard_keys (
		.clk      (clk_25_in_clk),                                            //                 clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),                      //               reset.reset_n
		.address  (keyboard_keys_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (keyboard_keys_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (keyboard_keys_export)                                      // external_connection.export
	);

	DE2_QSYS_modulation_selector modulation_selector (
		.clk        (clk_clk),                                                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                                  //               reset.reset_n
		.address    (modulation_selector_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~modulation_selector_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (modulation_selector_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (modulation_selector_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (modulation_selector_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (modulation_selector_export)                                        // external_connection.export
	);

	DE2_QSYS_mouse_pos mouse_pos (
		.clk      (clk_40_in_clk),                                        //                 clk.clk
		.reset_n  (~rst_controller_003_reset_out_reset),                  //               reset.reset_n
		.address  (mouse_pos_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (mouse_pos_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (mouse_pos_export)                                      // external_connection.export
	);

	DE2_QSYS_sdram sdram (
		.clk            (cpu_clk_for_sdram_clk),                                 //   clk.clk
		.reset_n        (~rst_controller_004_reset_out_reset),                   // reset.reset_n
		.az_addr        (sdram_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~sdram_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (sdram_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (sdram_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~sdram_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~sdram_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (sdram_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (sdram_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (sdram_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                                       //  wire.export
		.zs_ba          (sdram_wire_ba),                                         //      .export
		.zs_cas_n       (sdram_wire_cas_n),                                      //      .export
		.zs_cke         (sdram_wire_cke),                                        //      .export
		.zs_cs_n        (sdram_wire_cs_n),                                       //      .export
		.zs_dq          (sdram_wire_dq),                                         //      .export
		.zs_dqm         (sdram_wire_dqm),                                        //      .export
		.zs_ras_n       (sdram_wire_ras_n),                                      //      .export
		.zs_we_n        (sdram_wire_we_n)                                        //      .export
	);

	DE2_QSYS_signal_selector signal_selector (
		.clk        (clk_clk),                                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                              //               reset.reset_n
		.address    (signal_selector_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~signal_selector_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (signal_selector_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (signal_selector_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (signal_selector_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (signal_selector_export)                                        // external_connection.export
	);

	DE2_QSYS_sysid_qsys sysid_qsys (
		.clock    (clk_clk),                                                          //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                                  //         reset.reset_n
		.readdata (sysid_qsys_control_slave_translator_avalon_anti_slave_0_readdata), // control_slave.readdata
		.address  (sysid_qsys_control_slave_translator_avalon_anti_slave_0_address)   //              .address
	);

	DE2_QSYS_timer timer (
		.clk        (clk_clk),                                            //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    // reset.reset_n
		.address    (timer_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                            //   irq.irq
	);

	DE2_QSYS_vga vga (
		.alt_vip_itc_0_clocked_video_vid_clk       (vga_alt_vip_itc_0_clocked_video_vid_clk),                           //    alt_vip_itc_0_clocked_video.vid_clk
		.alt_vip_itc_0_clocked_video_vid_data      (vga_alt_vip_itc_0_clocked_video_vid_data),                          //                               .vid_data
		.alt_vip_itc_0_clocked_video_underflow     (vga_alt_vip_itc_0_clocked_video_underflow),                         //                               .underflow
		.alt_vip_itc_0_clocked_video_vid_datavalid (vga_alt_vip_itc_0_clocked_video_vid_datavalid),                     //                               .vid_datavalid
		.alt_vip_itc_0_clocked_video_vid_v_sync    (vga_alt_vip_itc_0_clocked_video_vid_v_sync),                        //                               .vid_v_sync
		.alt_vip_itc_0_clocked_video_vid_h_sync    (vga_alt_vip_itc_0_clocked_video_vid_h_sync),                        //                               .vid_h_sync
		.alt_vip_itc_0_clocked_video_vid_f         (vga_alt_vip_itc_0_clocked_video_vid_f),                             //                               .vid_f
		.alt_vip_itc_0_clocked_video_vid_h         (vga_alt_vip_itc_0_clocked_video_vid_h),                             //                               .vid_h
		.alt_vip_itc_0_clocked_video_vid_v         (vga_alt_vip_itc_0_clocked_video_vid_v),                             //                               .vid_v
		.alt_vip_vfr_0_interrupt_sender_irq        (irq_synchronizer_receiver_irq),                                     // alt_vip_vfr_0_interrupt_sender.irq
		.nios_clk_clk                              (cpu_clk_for_sdram_clk),                                             //                       nios_clk.clk
		.nios_clk_reset_reset_n                    (reset_reset_n),                                                     //                 nios_clk_reset.reset_n
		.to_nios_2_datamaster_address              (vga_to_nios_2_datamaster_translator_avalon_anti_slave_0_address),   //           to_nios_2_datamaster.address
		.to_nios_2_datamaster_write                (vga_to_nios_2_datamaster_translator_avalon_anti_slave_0_write),     //                               .write
		.to_nios_2_datamaster_writedata            (vga_to_nios_2_datamaster_translator_avalon_anti_slave_0_writedata), //                               .writedata
		.to_nios_2_datamaster_read                 (vga_to_nios_2_datamaster_translator_avalon_anti_slave_0_read),      //                               .read
		.to_nios_2_datamaster_readdata             (vga_to_nios_2_datamaster_translator_avalon_anti_slave_0_readdata),  //                               .readdata
		.to_sdram_address                          (vga_to_sdram_address),                                              //                       to_sdram.address
		.to_sdram_burstcount                       (vga_to_sdram_burstcount),                                           //                               .burstcount
		.to_sdram_readdata                         (vga_to_sdram_readdata),                                             //                               .readdata
		.to_sdram_read                             (vga_to_sdram_read),                                                 //                               .read
		.to_sdram_readdatavalid                    (vga_to_sdram_readdatavalid),                                        //                               .readdatavalid
		.to_sdram_waitrequest                      (vga_to_sdram_waitrequest)                                           //                               .waitrequest
	);

	DE2_QSYS_lfsr_clk_interrupt_gen lfsr_clk_interrupt_gen (
		.clk        (clk_clk),                                                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                                     //               reset.reset_n
		.address    (lfsr_clk_interrupt_gen_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~lfsr_clk_interrupt_gen_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (lfsr_clk_interrupt_gen_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (lfsr_clk_interrupt_gen_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (lfsr_clk_interrupt_gen_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (lfsr_clk_interrupt_gen_external_connection_export),                   // external_connection.export
		.irq        ()                                                                     //                 irq.irq
	);

	DE2_QSYS_lfsr_val lfsr_val (
		.clk      (clk_clk),                                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                     //               reset.reset_n
		.address  (lfsr_val_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (lfsr_val_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (lfsr_val_external_connection_export)                  // external_connection.export
	);

	DE2_QSYS_div_freq dds_increment (
		.clk        (clk_clk),                                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                            //               reset.reset_n
		.address    (dds_increment_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~dds_increment_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (dds_increment_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (dds_increment_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (dds_increment_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (dds_increment_external_connection_export)                    // external_connection.export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (25),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_data_master_translator (
		.clk                      (clk_clk),                                                            //                       clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                 //                     reset.reset
		.uav_address              (cpu_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (cpu_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (cpu_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (cpu_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (cpu_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (cpu_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (cpu_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (cpu_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (cpu_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (cpu_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (cpu_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (cpu_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (cpu_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (cpu_data_master_byteenable),                                         //                          .byteenable
		.av_read                  (cpu_data_master_read),                                               //                          .read
		.av_readdata              (cpu_data_master_readdata),                                           //                          .readdata
		.av_write                 (cpu_data_master_write),                                              //                          .write
		.av_writedata             (cpu_data_master_writedata),                                          //                          .writedata
		.av_debugaccess           (cpu_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount            (1'b1),                                                               //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                               //               (terminated)
		.av_begintransfer         (1'b0),                                                               //               (terminated)
		.av_chipselect            (1'b0),                                                               //               (terminated)
		.av_readdatavalid         (),                                                                   //               (terminated)
		.av_lock                  (1'b0),                                                               //               (terminated)
		.uav_clken                (),                                                                   //               (terminated)
		.av_clken                 (1'b1),                                                               //               (terminated)
		.uav_response             (2'b00),                                                              //               (terminated)
		.av_response              (),                                                                   //               (terminated)
		.uav_writeresponserequest (),                                                                   //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                               //               (terminated)
		.av_writeresponserequest  (1'b0),                                                               //               (terminated)
		.av_writeresponsevalid    ()                                                                    //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (6),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (8),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (1),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) vga_to_sdram_translator (
		.clk                      (cpu_clk_for_sdram_clk),                                           //                       clk.clk
		.reset                    (rst_controller_004_reset_out_reset),                              //                     reset.reset
		.uav_address              (vga_to_sdram_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (vga_to_sdram_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (vga_to_sdram_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (vga_to_sdram_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (vga_to_sdram_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (vga_to_sdram_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (vga_to_sdram_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (vga_to_sdram_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (vga_to_sdram_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (vga_to_sdram_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (vga_to_sdram_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (vga_to_sdram_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (vga_to_sdram_waitrequest),                                        //                          .waitrequest
		.av_burstcount            (vga_to_sdram_burstcount),                                         //                          .burstcount
		.av_read                  (vga_to_sdram_read),                                               //                          .read
		.av_readdata              (vga_to_sdram_readdata),                                           //                          .readdata
		.av_readdatavalid         (vga_to_sdram_readdatavalid),                                      //                          .readdatavalid
		.av_byteenable            (4'b1111),                                                         //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                            //               (terminated)
		.av_begintransfer         (1'b0),                                                            //               (terminated)
		.av_chipselect            (1'b0),                                                            //               (terminated)
		.av_write                 (1'b0),                                                            //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                            //               (terminated)
		.av_lock                  (1'b0),                                                            //               (terminated)
		.av_debugaccess           (1'b0),                                                            //               (terminated)
		.uav_clken                (),                                                                //               (terminated)
		.av_clken                 (1'b1),                                                            //               (terminated)
		.uav_response             (2'b00),                                                           //               (terminated)
		.av_response              (),                                                                //               (terminated)
		.uav_writeresponserequest (),                                                                //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                            //               (terminated)
		.av_writeresponserequest  (1'b0),                                                            //               (terminated)
		.av_writeresponsevalid    ()                                                                 //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (25),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_instruction_master_translator (
		.clk                      (clk_clk),                                                                   //                       clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                        //                     reset.reset
		.uav_address              (cpu_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (cpu_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (cpu_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (cpu_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (cpu_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (cpu_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (cpu_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (cpu_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (cpu_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (cpu_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (cpu_instruction_master_read),                                               //                          .read
		.av_readdata              (cpu_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (cpu_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount            (1'b1),                                                                      //               (terminated)
		.av_byteenable            (4'b1111),                                                                   //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                      //               (terminated)
		.av_begintransfer         (1'b0),                                                                      //               (terminated)
		.av_chipselect            (1'b0),                                                                      //               (terminated)
		.av_write                 (1'b0),                                                                      //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                      //               (terminated)
		.av_lock                  (1'b0),                                                                      //               (terminated)
		.av_debugaccess           (1'b0),                                                                      //               (terminated)
		.uav_clken                (),                                                                          //               (terminated)
		.av_clken                 (1'b1),                                                                      //               (terminated)
		.uav_response             (2'b00),                                                                     //               (terminated)
		.av_response              (),                                                                          //               (terminated)
		.uav_writeresponserequest (),                                                                          //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                      //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                      //               (terminated)
		.av_writeresponsevalid    ()                                                                           //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_avalon_jtag_slave_translator (
		.clk                      (clk_clk),                                                                                //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                         //                    reset.reset
		.uav_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                                       //              (terminated)
		.av_burstcount            (),                                                                                       //              (terminated)
		.av_byteenable            (),                                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                                       //              (terminated)
		.av_lock                  (),                                                                                       //              (terminated)
		.av_clken                 (),                                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                                   //              (terminated)
		.av_debugaccess           (),                                                                                       //              (terminated)
		.av_outputenable          (),                                                                                       //              (terminated)
		.uav_response             (),                                                                                       //              (terminated)
		.av_response              (2'b00),                                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sysid_qsys_control_slave_translator (
		.clk                      (clk_clk),                                                                             //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                      //                    reset.reset
		.uav_address              (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sysid_qsys_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (sysid_qsys_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                                    //              (terminated)
		.av_read                  (),                                                                                    //              (terminated)
		.av_writedata             (),                                                                                    //              (terminated)
		.av_begintransfer         (),                                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                                    //              (terminated)
		.av_burstcount            (),                                                                                    //              (terminated)
		.av_byteenable            (),                                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                                //              (terminated)
		.av_writebyteenable       (),                                                                                    //              (terminated)
		.av_lock                  (),                                                                                    //              (terminated)
		.av_chipselect            (),                                                                                    //              (terminated)
		.av_clken                 (),                                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                                //              (terminated)
		.av_debugaccess           (),                                                                                    //              (terminated)
		.av_outputenable          (),                                                                                    //              (terminated)
		.uav_response             (),                                                                                    //              (terminated)
		.av_response              (2'b00),                                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) audio_data_fregen_s1_translator (
		.clk                      (clk_clk),                                                                         //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                  //                    reset.reset
		.uav_address              (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (audio_data_fregen_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (audio_data_fregen_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (audio_data_fregen_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (audio_data_fregen_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (audio_data_fregen_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                                //              (terminated)
		.av_begintransfer         (),                                                                                //              (terminated)
		.av_beginbursttransfer    (),                                                                                //              (terminated)
		.av_burstcount            (),                                                                                //              (terminated)
		.av_byteenable            (),                                                                                //              (terminated)
		.av_readdatavalid         (1'b0),                                                                            //              (terminated)
		.av_waitrequest           (1'b0),                                                                            //              (terminated)
		.av_writebyteenable       (),                                                                                //              (terminated)
		.av_lock                  (),                                                                                //              (terminated)
		.av_clken                 (),                                                                                //              (terminated)
		.uav_clken                (1'b0),                                                                            //              (terminated)
		.av_debugaccess           (),                                                                                //              (terminated)
		.av_outputenable          (),                                                                                //              (terminated)
		.uav_response             (),                                                                                //              (terminated)
		.av_response              (2'b00),                                                                           //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                            //              (terminated)
		.uav_writeresponsevalid   (),                                                                                //              (terminated)
		.av_writeresponserequest  (),                                                                                //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) audio_empty_s1_translator (
		.clk                      (clk_clk),                                                                   //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                            //                    reset.reset
		.uav_address              (audio_empty_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (audio_empty_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (audio_empty_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (audio_empty_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (audio_empty_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (audio_empty_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (audio_empty_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (audio_empty_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (audio_empty_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (audio_empty_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (audio_empty_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (audio_empty_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (audio_empty_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                          //              (terminated)
		.av_read                  (),                                                                          //              (terminated)
		.av_writedata             (),                                                                          //              (terminated)
		.av_begintransfer         (),                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                          //              (terminated)
		.av_burstcount            (),                                                                          //              (terminated)
		.av_byteenable            (),                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                      //              (terminated)
		.av_waitrequest           (1'b0),                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                          //              (terminated)
		.av_lock                  (),                                                                          //              (terminated)
		.av_chipselect            (),                                                                          //              (terminated)
		.av_clken                 (),                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                      //              (terminated)
		.av_debugaccess           (),                                                                          //              (terminated)
		.av_outputenable          (),                                                                          //              (terminated)
		.uav_response             (),                                                                          //              (terminated)
		.av_response              (2'b00),                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) audio_fifo_full_s1_translator (
		.clk                      (clk_clk),                                                                       //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                //                    reset.reset
		.uav_address              (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (audio_fifo_full_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (audio_fifo_full_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                              //              (terminated)
		.av_read                  (),                                                                              //              (terminated)
		.av_writedata             (),                                                                              //              (terminated)
		.av_begintransfer         (),                                                                              //              (terminated)
		.av_beginbursttransfer    (),                                                                              //              (terminated)
		.av_burstcount            (),                                                                              //              (terminated)
		.av_byteenable            (),                                                                              //              (terminated)
		.av_readdatavalid         (1'b0),                                                                          //              (terminated)
		.av_waitrequest           (1'b0),                                                                          //              (terminated)
		.av_writebyteenable       (),                                                                              //              (terminated)
		.av_lock                  (),                                                                              //              (terminated)
		.av_chipselect            (),                                                                              //              (terminated)
		.av_clken                 (),                                                                              //              (terminated)
		.uav_clken                (1'b0),                                                                          //              (terminated)
		.av_debugaccess           (),                                                                              //              (terminated)
		.av_outputenable          (),                                                                              //              (terminated)
		.uav_response             (),                                                                              //              (terminated)
		.av_response              (2'b00),                                                                         //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                          //              (terminated)
		.uav_writeresponsevalid   (),                                                                              //              (terminated)
		.av_writeresponserequest  (),                                                                              //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) audio_fifo_used_s1_translator (
		.clk                      (clk_clk),                                                                       //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                //                    reset.reset
		.uav_address              (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (audio_fifo_used_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (audio_fifo_used_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                              //              (terminated)
		.av_read                  (),                                                                              //              (terminated)
		.av_writedata             (),                                                                              //              (terminated)
		.av_begintransfer         (),                                                                              //              (terminated)
		.av_beginbursttransfer    (),                                                                              //              (terminated)
		.av_burstcount            (),                                                                              //              (terminated)
		.av_byteenable            (),                                                                              //              (terminated)
		.av_readdatavalid         (1'b0),                                                                          //              (terminated)
		.av_waitrequest           (1'b0),                                                                          //              (terminated)
		.av_writebyteenable       (),                                                                              //              (terminated)
		.av_lock                  (),                                                                              //              (terminated)
		.av_chipselect            (),                                                                              //              (terminated)
		.av_clken                 (),                                                                              //              (terminated)
		.uav_clken                (1'b0),                                                                          //              (terminated)
		.av_debugaccess           (),                                                                              //              (terminated)
		.av_outputenable          (),                                                                              //              (terminated)
		.uav_response             (),                                                                              //              (terminated)
		.av_response              (2'b00),                                                                         //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                          //              (terminated)
		.uav_writeresponsevalid   (),                                                                              //              (terminated)
		.av_writeresponserequest  (),                                                                              //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_jtag_debug_module_translator (
		.clk                      (clk_clk),                                                                          //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                               //                    reset.reset
		.uav_address              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (cpu_jtag_debug_module_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                 //              (terminated)
		.av_beginbursttransfer    (),                                                                                 //              (terminated)
		.av_burstcount            (),                                                                                 //              (terminated)
		.av_readdatavalid         (1'b0),                                                                             //              (terminated)
		.av_writebyteenable       (),                                                                                 //              (terminated)
		.av_lock                  (),                                                                                 //              (terminated)
		.av_chipselect            (),                                                                                 //              (terminated)
		.av_clken                 (),                                                                                 //              (terminated)
		.uav_clken                (1'b0),                                                                             //              (terminated)
		.av_outputenable          (),                                                                                 //              (terminated)
		.uav_response             (),                                                                                 //              (terminated)
		.av_response              (2'b00),                                                                            //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                             //              (terminated)
		.uav_writeresponsevalid   (),                                                                                 //              (terminated)
		.av_writeresponserequest  (),                                                                                 //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) audio_out_data_audio_s1_translator (
		.clk                      (clk_clk),                                                                            //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                     //                    reset.reset
		.uav_address              (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (audio_out_data_audio_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (audio_out_data_audio_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (audio_out_data_audio_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (audio_out_data_audio_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (audio_out_data_audio_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                                   //              (terminated)
		.av_begintransfer         (),                                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                                   //              (terminated)
		.av_burstcount            (),                                                                                   //              (terminated)
		.av_byteenable            (),                                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                                               //              (terminated)
		.av_writebyteenable       (),                                                                                   //              (terminated)
		.av_lock                  (),                                                                                   //              (terminated)
		.av_clken                 (),                                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                                               //              (terminated)
		.av_debugaccess           (),                                                                                   //              (terminated)
		.av_outputenable          (),                                                                                   //              (terminated)
		.uav_response             (),                                                                                   //              (terminated)
		.av_response              (2'b00),                                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) audio_out_pause_s1_translator (
		.clk                      (clk_clk),                                                                       //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                //                    reset.reset
		.uav_address              (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (audio_out_pause_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (audio_out_pause_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (audio_out_pause_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (audio_out_pause_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (audio_out_pause_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                              //              (terminated)
		.av_begintransfer         (),                                                                              //              (terminated)
		.av_beginbursttransfer    (),                                                                              //              (terminated)
		.av_burstcount            (),                                                                              //              (terminated)
		.av_byteenable            (),                                                                              //              (terminated)
		.av_readdatavalid         (1'b0),                                                                          //              (terminated)
		.av_waitrequest           (1'b0),                                                                          //              (terminated)
		.av_writebyteenable       (),                                                                              //              (terminated)
		.av_lock                  (),                                                                              //              (terminated)
		.av_clken                 (),                                                                              //              (terminated)
		.uav_clken                (1'b0),                                                                          //              (terminated)
		.av_debugaccess           (),                                                                              //              (terminated)
		.av_outputenable          (),                                                                              //              (terminated)
		.uav_response             (),                                                                              //              (terminated)
		.av_response              (2'b00),                                                                         //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                          //              (terminated)
		.uav_writeresponsevalid   (),                                                                              //              (terminated)
		.av_writeresponserequest  (),                                                                              //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) audio_out_stop_s1_translator (
		.clk                      (clk_clk),                                                                      //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                               //                    reset.reset
		.uav_address              (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (audio_out_stop_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (audio_out_stop_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (audio_out_stop_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (audio_out_stop_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (audio_out_stop_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                             //              (terminated)
		.av_begintransfer         (),                                                                             //              (terminated)
		.av_beginbursttransfer    (),                                                                             //              (terminated)
		.av_burstcount            (),                                                                             //              (terminated)
		.av_byteenable            (),                                                                             //              (terminated)
		.av_readdatavalid         (1'b0),                                                                         //              (terminated)
		.av_waitrequest           (1'b0),                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                             //              (terminated)
		.av_lock                  (),                                                                             //              (terminated)
		.av_clken                 (),                                                                             //              (terminated)
		.uav_clken                (1'b0),                                                                         //              (terminated)
		.av_debugaccess           (),                                                                             //              (terminated)
		.av_outputenable          (),                                                                             //              (terminated)
		.uav_response             (),                                                                             //              (terminated)
		.av_response              (2'b00),                                                                        //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                         //              (terminated)
		.uav_writeresponsevalid   (),                                                                             //              (terminated)
		.av_writeresponserequest  (),                                                                             //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_s1_translator (
		.clk                      (clk_clk),                                                             //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                      //                    reset.reset
		.uav_address              (timer_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (timer_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (timer_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (timer_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (timer_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (timer_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (timer_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                    //              (terminated)
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_byteenable            (),                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) key_s1_translator (
		.clk                      (clk_clk),                                                           //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                    //                    reset.reset
		.uav_address              (key_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (key_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (key_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (key_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (key_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (key_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (key_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (key_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (key_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (key_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (key_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (key_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (key_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (key_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (key_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (key_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                  //              (terminated)
		.av_begintransfer         (),                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                  //              (terminated)
		.av_burstcount            (),                                                                  //              (terminated)
		.av_byteenable            (),                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                              //              (terminated)
		.av_waitrequest           (1'b0),                                                              //              (terminated)
		.av_writebyteenable       (),                                                                  //              (terminated)
		.av_lock                  (),                                                                  //              (terminated)
		.av_clken                 (),                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                              //              (terminated)
		.av_debugaccess           (),                                                                  //              (terminated)
		.av_outputenable          (),                                                                  //              (terminated)
		.uav_response             (),                                                                  //              (terminated)
		.av_response              (2'b00),                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) signal_selector_s1_translator (
		.clk                      (clk_clk),                                                                       //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                //                    reset.reset
		.uav_address              (signal_selector_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (signal_selector_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (signal_selector_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (signal_selector_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (signal_selector_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (signal_selector_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (signal_selector_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (signal_selector_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (signal_selector_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (signal_selector_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (signal_selector_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (signal_selector_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (signal_selector_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (signal_selector_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (signal_selector_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (signal_selector_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                              //              (terminated)
		.av_begintransfer         (),                                                                              //              (terminated)
		.av_beginbursttransfer    (),                                                                              //              (terminated)
		.av_burstcount            (),                                                                              //              (terminated)
		.av_byteenable            (),                                                                              //              (terminated)
		.av_readdatavalid         (1'b0),                                                                          //              (terminated)
		.av_waitrequest           (1'b0),                                                                          //              (terminated)
		.av_writebyteenable       (),                                                                              //              (terminated)
		.av_lock                  (),                                                                              //              (terminated)
		.av_clken                 (),                                                                              //              (terminated)
		.uav_clken                (1'b0),                                                                          //              (terminated)
		.av_debugaccess           (),                                                                              //              (terminated)
		.av_outputenable          (),                                                                              //              (terminated)
		.uav_response             (),                                                                              //              (terminated)
		.av_response              (2'b00),                                                                         //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                          //              (terminated)
		.uav_writeresponsevalid   (),                                                                              //              (terminated)
		.av_writeresponserequest  (),                                                                              //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) modulation_selector_s1_translator (
		.clk                      (clk_clk),                                                                           //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                    //                    reset.reset
		.uav_address              (modulation_selector_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (modulation_selector_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (modulation_selector_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (modulation_selector_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (modulation_selector_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (modulation_selector_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (modulation_selector_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (modulation_selector_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (modulation_selector_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (modulation_selector_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (modulation_selector_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (modulation_selector_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (modulation_selector_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (modulation_selector_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (modulation_selector_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (modulation_selector_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                                  //              (terminated)
		.av_begintransfer         (),                                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                                  //              (terminated)
		.av_burstcount            (),                                                                                  //              (terminated)
		.av_byteenable            (),                                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                                              //              (terminated)
		.av_waitrequest           (1'b0),                                                                              //              (terminated)
		.av_writebyteenable       (),                                                                                  //              (terminated)
		.av_lock                  (),                                                                                  //              (terminated)
		.av_clken                 (),                                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                                              //              (terminated)
		.av_debugaccess           (),                                                                                  //              (terminated)
		.av_outputenable          (),                                                                                  //              (terminated)
		.uav_response             (),                                                                                  //              (terminated)
		.av_response              (2'b00),                                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) keyboard_keys_s1_translator (
		.clk                      (clk_25_in_clk),                                                               //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                          //                    reset.reset
		.uav_address              (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (keyboard_keys_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (keyboard_keys_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                            //              (terminated)
		.av_read                  (),                                                                            //              (terminated)
		.av_writedata             (),                                                                            //              (terminated)
		.av_begintransfer         (),                                                                            //              (terminated)
		.av_beginbursttransfer    (),                                                                            //              (terminated)
		.av_burstcount            (),                                                                            //              (terminated)
		.av_byteenable            (),                                                                            //              (terminated)
		.av_readdatavalid         (1'b0),                                                                        //              (terminated)
		.av_waitrequest           (1'b0),                                                                        //              (terminated)
		.av_writebyteenable       (),                                                                            //              (terminated)
		.av_lock                  (),                                                                            //              (terminated)
		.av_chipselect            (),                                                                            //              (terminated)
		.av_clken                 (),                                                                            //              (terminated)
		.uav_clken                (1'b0),                                                                        //              (terminated)
		.av_debugaccess           (),                                                                            //              (terminated)
		.av_outputenable          (),                                                                            //              (terminated)
		.uav_response             (),                                                                            //              (terminated)
		.av_response              (2'b00),                                                                       //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                        //              (terminated)
		.uav_writeresponsevalid   (),                                                                            //              (terminated)
		.av_writeresponserequest  (),                                                                            //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) mouse_pos_s1_translator (
		.clk                      (clk_40_in_clk),                                                           //                      clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                      //                    reset.reset
		.uav_address              (mouse_pos_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (mouse_pos_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (mouse_pos_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (mouse_pos_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (mouse_pos_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (mouse_pos_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (mouse_pos_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (mouse_pos_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (mouse_pos_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (mouse_pos_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (mouse_pos_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (mouse_pos_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (mouse_pos_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                        //              (terminated)
		.av_read                  (),                                                                        //              (terminated)
		.av_writedata             (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_chipselect            (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) div_freq_s1_translator (
		.clk                      (clk_clk),                                                                //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                         //                    reset.reset
		.uav_address              (div_freq_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (div_freq_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (div_freq_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (div_freq_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (div_freq_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (div_freq_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (div_freq_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (div_freq_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (div_freq_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (div_freq_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (div_freq_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (div_freq_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (div_freq_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (div_freq_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (div_freq_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (div_freq_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                       //              (terminated)
		.av_begintransfer         (),                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                       //              (terminated)
		.av_burstcount            (),                                                                       //              (terminated)
		.av_byteenable            (),                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                   //              (terminated)
		.av_waitrequest           (1'b0),                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                       //              (terminated)
		.av_lock                  (),                                                                       //              (terminated)
		.av_clken                 (),                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                   //              (terminated)
		.av_debugaccess           (),                                                                       //              (terminated)
		.av_outputenable          (),                                                                       //              (terminated)
		.uav_response             (),                                                                       //              (terminated)
		.av_response              (2'b00),                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) audio_sel_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                          //                    reset.reset
		.uav_address              (audio_sel_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (audio_sel_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (audio_sel_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (audio_sel_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (audio_sel_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (audio_sel_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (audio_sel_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (audio_sel_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (audio_sel_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (audio_sel_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (audio_sel_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (audio_sel_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (audio_sel_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (audio_sel_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (audio_sel_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (audio_sel_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (5),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) vga_to_nios_2_datamaster_translator (
		.clk                      (cpu_clk_for_sdram_clk),                                                               //                      clk.clk
		.reset                    (rst_controller_004_reset_out_reset),                                                  //                    reset.reset
		.uav_address              (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (vga_to_nios_2_datamaster_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (vga_to_nios_2_datamaster_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (vga_to_nios_2_datamaster_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (vga_to_nios_2_datamaster_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (vga_to_nios_2_datamaster_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (),                                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                                    //              (terminated)
		.av_burstcount            (),                                                                                    //              (terminated)
		.av_byteenable            (),                                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                                //              (terminated)
		.av_writebyteenable       (),                                                                                    //              (terminated)
		.av_lock                  (),                                                                                    //              (terminated)
		.av_chipselect            (),                                                                                    //              (terminated)
		.av_clken                 (),                                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                                //              (terminated)
		.av_debugaccess           (),                                                                                    //              (terminated)
		.av_outputenable          (),                                                                                    //              (terminated)
		.uav_response             (),                                                                                    //              (terminated)
		.av_response              (2'b00),                                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) audio_wrclk_s1_translator (
		.clk                      (clk_clk),                                                                   //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                            //                    reset.reset
		.uav_address              (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (audio_wrclk_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (audio_wrclk_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (audio_wrclk_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (audio_wrclk_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (audio_wrclk_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                          //              (terminated)
		.av_begintransfer         (),                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                          //              (terminated)
		.av_burstcount            (),                                                                          //              (terminated)
		.av_byteenable            (),                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                      //              (terminated)
		.av_waitrequest           (1'b0),                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                          //              (terminated)
		.av_lock                  (),                                                                          //              (terminated)
		.av_clken                 (),                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                      //              (terminated)
		.av_debugaccess           (),                                                                          //              (terminated)
		.av_outputenable          (),                                                                          //              (terminated)
		.uav_response             (),                                                                          //              (terminated)
		.av_response              (2'b00),                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) audio_wrreq_s1_translator (
		.clk                      (clk_clk),                                                                   //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                            //                    reset.reset
		.uav_address              (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (audio_wrreq_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (audio_wrreq_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (audio_wrreq_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (audio_wrreq_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (audio_wrreq_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                          //              (terminated)
		.av_begintransfer         (),                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                          //              (terminated)
		.av_burstcount            (),                                                                          //              (terminated)
		.av_byteenable            (),                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                      //              (terminated)
		.av_waitrequest           (1'b0),                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                          //              (terminated)
		.av_lock                  (),                                                                          //              (terminated)
		.av_clken                 (),                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                      //              (terminated)
		.av_debugaccess           (),                                                                          //              (terminated)
		.av_outputenable          (),                                                                          //              (terminated)
		.uav_response             (),                                                                          //              (terminated)
		.av_response              (2'b00),                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (22),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sdram_s1_translator (
		.clk                      (cpu_clk_for_sdram_clk),                                               //                      clk.clk
		.reset                    (rst_controller_004_reset_out_reset),                                  //                    reset.reset
		.uav_address              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sdram_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (sdram_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (sdram_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (sdram_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (sdram_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (sdram_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (sdram_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (sdram_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (sdram_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) lfsr_clk_interrupt_gen_s1_translator (
		.clk                      (clk_clk),                                                                              //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                       //                    reset.reset
		.uav_address              (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (lfsr_clk_interrupt_gen_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (lfsr_clk_interrupt_gen_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (lfsr_clk_interrupt_gen_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (lfsr_clk_interrupt_gen_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (lfsr_clk_interrupt_gen_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                                     //              (terminated)
		.av_begintransfer         (),                                                                                     //              (terminated)
		.av_beginbursttransfer    (),                                                                                     //              (terminated)
		.av_burstcount            (),                                                                                     //              (terminated)
		.av_byteenable            (),                                                                                     //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                 //              (terminated)
		.av_waitrequest           (1'b0),                                                                                 //              (terminated)
		.av_writebyteenable       (),                                                                                     //              (terminated)
		.av_lock                  (),                                                                                     //              (terminated)
		.av_clken                 (),                                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                                 //              (terminated)
		.av_debugaccess           (),                                                                                     //              (terminated)
		.av_outputenable          (),                                                                                     //              (terminated)
		.uav_response             (),                                                                                     //              (terminated)
		.av_response              (2'b00),                                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) lfsr_val_s1_translator (
		.clk                      (clk_clk),                                                                //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                         //                    reset.reset
		.uav_address              (lfsr_val_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (lfsr_val_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (lfsr_val_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (lfsr_val_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (lfsr_val_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (lfsr_val_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (lfsr_val_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (lfsr_val_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (lfsr_val_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (lfsr_val_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (lfsr_val_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (lfsr_val_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (lfsr_val_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                       //              (terminated)
		.av_read                  (),                                                                       //              (terminated)
		.av_writedata             (),                                                                       //              (terminated)
		.av_begintransfer         (),                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                       //              (terminated)
		.av_burstcount            (),                                                                       //              (terminated)
		.av_byteenable            (),                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                   //              (terminated)
		.av_waitrequest           (1'b0),                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                       //              (terminated)
		.av_lock                  (),                                                                       //              (terminated)
		.av_chipselect            (),                                                                       //              (terminated)
		.av_clken                 (),                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                   //              (terminated)
		.av_debugaccess           (),                                                                       //              (terminated)
		.av_outputenable          (),                                                                       //              (terminated)
		.uav_response             (),                                                                       //              (terminated)
		.av_response              (2'b00),                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) dds_increment_s1_translator (
		.clk                      (clk_clk),                                                                     //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                              //                    reset.reset
		.uav_address              (dds_increment_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (dds_increment_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (dds_increment_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (dds_increment_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (dds_increment_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (dds_increment_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (dds_increment_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (dds_increment_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (dds_increment_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (dds_increment_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (dds_increment_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (dds_increment_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (dds_increment_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (dds_increment_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (dds_increment_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (dds_increment_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                            //              (terminated)
		.av_begintransfer         (),                                                                            //              (terminated)
		.av_beginbursttransfer    (),                                                                            //              (terminated)
		.av_burstcount            (),                                                                            //              (terminated)
		.av_byteenable            (),                                                                            //              (terminated)
		.av_readdatavalid         (1'b0),                                                                        //              (terminated)
		.av_waitrequest           (1'b0),                                                                        //              (terminated)
		.av_writebyteenable       (),                                                                            //              (terminated)
		.av_lock                  (),                                                                            //              (terminated)
		.av_clken                 (),                                                                            //              (terminated)
		.uav_clken                (1'b0),                                                                        //              (terminated)
		.av_debugaccess           (),                                                                            //              (terminated)
		.av_outputenable          (),                                                                            //              (terminated)
		.uav_response             (),                                                                            //              (terminated)
		.av_response              (2'b00),                                                                       //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                        //              (terminated)
		.uav_writeresponsevalid   (),                                                                            //              (terminated)
		.av_writeresponserequest  (),                                                                            //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                         //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (107),
		.PKT_PROTECTION_L          (105),
		.PKT_BEGIN_BURST           (92),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.PKT_BURST_TYPE_H          (89),
		.PKT_BURST_TYPE_L          (88),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (103),
		.PKT_DEST_ID_L             (99),
		.PKT_THREAD_ID_H           (104),
		.PKT_THREAD_ID_L           (104),
		.PKT_CACHE_H               (111),
		.PKT_CACHE_L               (108),
		.PKT_DATA_SIDEBAND_H       (91),
		.PKT_DATA_SIDEBAND_L       (91),
		.PKT_QOS_H                 (93),
		.PKT_QOS_L                 (93),
		.PKT_ADDR_SIDEBAND_H       (90),
		.PKT_ADDR_SIDEBAND_L       (90),
		.PKT_RESPONSE_STATUS_H     (113),
		.PKT_RESPONSE_STATUS_L     (112),
		.ST_DATA_W                 (114),
		.ST_CHANNEL_W              (25),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cpu_data_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                     //       clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.av_address              (cpu_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (cpu_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (cpu_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (cpu_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (cpu_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (cpu_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (cpu_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (cpu_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (cpu_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (cpu_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (cpu_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_src_valid),                                                      //        rp.valid
		.rp_data                 (rsp_xbar_mux_src_data),                                                       //          .data
		.rp_channel              (rsp_xbar_mux_src_channel),                                                    //          .channel
		.rp_startofpacket        (rsp_xbar_mux_src_startofpacket),                                              //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_src_endofpacket),                                                //          .endofpacket
		.rp_ready                (rsp_xbar_mux_src_ready),                                                      //          .ready
		.av_response             (),                                                                            // (terminated)
		.av_writeresponserequest (1'b0),                                                                        // (terminated)
		.av_writeresponsevalid   ()                                                                             // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (107),
		.PKT_PROTECTION_L          (105),
		.PKT_BEGIN_BURST           (92),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.PKT_BURST_TYPE_H          (89),
		.PKT_BURST_TYPE_L          (88),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (103),
		.PKT_DEST_ID_L             (99),
		.PKT_THREAD_ID_H           (104),
		.PKT_THREAD_ID_L           (104),
		.PKT_CACHE_H               (111),
		.PKT_CACHE_L               (108),
		.PKT_DATA_SIDEBAND_H       (91),
		.PKT_DATA_SIDEBAND_L       (91),
		.PKT_QOS_H                 (93),
		.PKT_QOS_L                 (93),
		.PKT_ADDR_SIDEBAND_H       (90),
		.PKT_ADDR_SIDEBAND_L       (90),
		.PKT_RESPONSE_STATUS_H     (113),
		.PKT_RESPONSE_STATUS_L     (112),
		.ST_DATA_W                 (114),
		.ST_CHANNEL_W              (25),
		.AV_BURSTCOUNT_W           (8),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (2),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) vga_to_sdram_translator_avalon_universal_master_0_agent (
		.clk                     (cpu_clk_for_sdram_clk),                                                    //       clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                       // clk_reset.reset
		.av_address              (vga_to_sdram_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (vga_to_sdram_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (vga_to_sdram_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (vga_to_sdram_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (vga_to_sdram_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (vga_to_sdram_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (vga_to_sdram_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (vga_to_sdram_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (vga_to_sdram_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (vga_to_sdram_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (vga_to_sdram_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (vga_to_sdram_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (vga_to_sdram_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (vga_to_sdram_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (vga_to_sdram_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (vga_to_sdram_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_demux_021_src1_valid),                                            //        rp.valid
		.rp_data                 (rsp_xbar_demux_021_src1_data),                                             //          .data
		.rp_channel              (rsp_xbar_demux_021_src1_channel),                                          //          .channel
		.rp_startofpacket        (rsp_xbar_demux_021_src1_startofpacket),                                    //          .startofpacket
		.rp_endofpacket          (rsp_xbar_demux_021_src1_endofpacket),                                      //          .endofpacket
		.rp_ready                (rsp_xbar_demux_021_src1_ready),                                            //          .ready
		.av_response             (),                                                                         // (terminated)
		.av_writeresponserequest (1'b0),                                                                     // (terminated)
		.av_writeresponsevalid   ()                                                                          // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (107),
		.PKT_PROTECTION_L          (105),
		.PKT_BEGIN_BURST           (92),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.PKT_BURST_TYPE_H          (89),
		.PKT_BURST_TYPE_L          (88),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (103),
		.PKT_DEST_ID_L             (99),
		.PKT_THREAD_ID_H           (104),
		.PKT_THREAD_ID_L           (104),
		.PKT_CACHE_H               (111),
		.PKT_CACHE_L               (108),
		.PKT_DATA_SIDEBAND_H       (91),
		.PKT_DATA_SIDEBAND_L       (91),
		.PKT_QOS_H                 (93),
		.PKT_QOS_L                 (93),
		.PKT_ADDR_SIDEBAND_H       (90),
		.PKT_ADDR_SIDEBAND_L       (90),
		.PKT_RESPONSE_STATUS_H     (113),
		.PKT_RESPONSE_STATUS_L     (112),
		.ST_DATA_W                 (114),
		.ST_CHANNEL_W              (25),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cpu_instruction_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                            //       clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.av_address              (cpu_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (cpu_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (cpu_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (cpu_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (cpu_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (cpu_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (cpu_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (cpu_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_rsp_src_valid),                                                              //        rp.valid
		.rp_data                 (limiter_rsp_src_data),                                                               //          .data
		.rp_channel              (limiter_rsp_src_channel),                                                            //          .channel
		.rp_startofpacket        (limiter_rsp_src_startofpacket),                                                      //          .startofpacket
		.rp_endofpacket          (limiter_rsp_src_endofpacket),                                                        //          .endofpacket
		.rp_ready                (limiter_rsp_src_ready),                                                              //          .ready
		.av_response             (),                                                                                   // (terminated)
		.av_writeresponserequest (1'b0),                                                                               // (terminated)
		.av_writeresponsevalid   ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (92),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (103),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (107),
		.PKT_PROTECTION_L          (105),
		.PKT_RESPONSE_STATUS_H     (113),
		.PKT_RESPONSE_STATUS_L     (112),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.ST_CHANNEL_W              (25),
		.ST_DATA_W                 (114),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                   //       clk_reset.reset
		.m0_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_source0_ready),                                                                     //              cp.ready
		.cp_valid                (agent_pipeline_source0_valid),                                                                     //                .valid
		.cp_data                 (agent_pipeline_source0_data),                                                                      //                .data
		.cp_startofpacket        (agent_pipeline_source0_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (agent_pipeline_source0_endofpacket),                                                               //                .endofpacket
		.cp_channel              (agent_pipeline_source0_channel),                                                                   //                .channel
		.rf_sink_ready           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (115),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                   // clk_reset.reset
		.in_data           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                             // clk_reset.reset
		.in_data           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_startofpacket  (1'b0),                                                                                       // (terminated)
		.in_endofpacket    (1'b0),                                                                                       // (terminated)
		.out_startofpacket (),                                                                                           // (terminated)
		.out_endofpacket   (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (92),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (103),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (107),
		.PKT_PROTECTION_L          (105),
		.PKT_RESPONSE_STATUS_H     (113),
		.PKT_RESPONSE_STATUS_L     (112),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.ST_CHANNEL_W              (25),
		.ST_DATA_W                 (114),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                       //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                //       clk_reset.reset
		.m0_address              (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_002_source0_ready),                                                              //              cp.ready
		.cp_valid                (agent_pipeline_002_source0_valid),                                                              //                .valid
		.cp_data                 (agent_pipeline_002_source0_data),                                                               //                .data
		.cp_startofpacket        (agent_pipeline_002_source0_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (agent_pipeline_002_source0_endofpacket),                                                        //                .endofpacket
		.cp_channel              (agent_pipeline_002_source0_channel),                                                            //                .channel
		.rf_sink_ready           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (115),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                // clk_reset.reset
		.in_data           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                          // (terminated)
		.csr_readdata      (),                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                          // (terminated)
		.almost_full_data  (),                                                                                              // (terminated)
		.almost_empty_data (),                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                          // (terminated)
		.out_empty         (),                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                          // (terminated)
		.out_error         (),                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                          // (terminated)
		.out_channel       ()                                                                                               // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_startofpacket  (1'b0),                                                                                    // (terminated)
		.in_endofpacket    (1'b0),                                                                                    // (terminated)
		.out_startofpacket (),                                                                                        // (terminated)
		.out_endofpacket   (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (92),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (103),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (107),
		.PKT_PROTECTION_L          (105),
		.PKT_RESPONSE_STATUS_H     (113),
		.PKT_RESPONSE_STATUS_L     (112),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.ST_CHANNEL_W              (25),
		.ST_DATA_W                 (114),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) audio_data_fregen_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                   //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                            //       clk_reset.reset
		.m0_address              (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_004_source0_ready),                                                          //              cp.ready
		.cp_valid                (agent_pipeline_004_source0_valid),                                                          //                .valid
		.cp_data                 (agent_pipeline_004_source0_data),                                                           //                .data
		.cp_startofpacket        (agent_pipeline_004_source0_startofpacket),                                                  //                .startofpacket
		.cp_endofpacket          (agent_pipeline_004_source0_endofpacket),                                                    //                .endofpacket
		.cp_channel              (agent_pipeline_004_source0_channel),                                                        //                .channel
		.rf_sink_ready           (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                     //     (terminated)
		.m0_writeresponserequest (),                                                                                          //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                       //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (115),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                   //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.in_data           (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                      // clk_reset.reset
		.in_data           (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_startofpacket  (1'b0),                                                                                // (terminated)
		.in_endofpacket    (1'b0),                                                                                // (terminated)
		.out_startofpacket (),                                                                                    // (terminated)
		.out_endofpacket   (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (92),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (103),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (107),
		.PKT_PROTECTION_L          (105),
		.PKT_RESPONSE_STATUS_H     (113),
		.PKT_RESPONSE_STATUS_L     (112),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.ST_CHANNEL_W              (25),
		.ST_DATA_W                 (114),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) audio_empty_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                             //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                      //       clk_reset.reset
		.m0_address              (audio_empty_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (audio_empty_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (audio_empty_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (audio_empty_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (audio_empty_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (audio_empty_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (audio_empty_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (audio_empty_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (audio_empty_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (audio_empty_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (audio_empty_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (audio_empty_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (audio_empty_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (audio_empty_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (audio_empty_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (audio_empty_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_006_source0_ready),                                                    //              cp.ready
		.cp_valid                (agent_pipeline_006_source0_valid),                                                    //                .valid
		.cp_data                 (agent_pipeline_006_source0_data),                                                     //                .data
		.cp_startofpacket        (agent_pipeline_006_source0_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (agent_pipeline_006_source0_endofpacket),                                              //                .endofpacket
		.cp_channel              (agent_pipeline_006_source0_channel),                                                  //                .channel
		.rf_sink_ready           (audio_empty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (audio_empty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (audio_empty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (audio_empty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (audio_empty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (audio_empty_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (audio_empty_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (audio_empty_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (audio_empty_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (audio_empty_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (audio_empty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (audio_empty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (audio_empty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (audio_empty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (audio_empty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (audio_empty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (115),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_empty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                      // clk_reset.reset
		.in_data           (audio_empty_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (audio_empty_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (audio_empty_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (audio_empty_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (audio_empty_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (audio_empty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (audio_empty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (audio_empty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (audio_empty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (audio_empty_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_empty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.in_data           (audio_empty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (audio_empty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (audio_empty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (audio_empty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (audio_empty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (audio_empty_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_startofpacket  (1'b0),                                                                          // (terminated)
		.in_endofpacket    (1'b0),                                                                          // (terminated)
		.out_startofpacket (),                                                                              // (terminated)
		.out_endofpacket   (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (92),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (103),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (107),
		.PKT_PROTECTION_L          (105),
		.PKT_RESPONSE_STATUS_H     (113),
		.PKT_RESPONSE_STATUS_L     (112),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.ST_CHANNEL_W              (25),
		.ST_DATA_W                 (114),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) audio_fifo_full_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                          //       clk_reset.reset
		.m0_address              (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_008_source0_ready),                                                        //              cp.ready
		.cp_valid                (agent_pipeline_008_source0_valid),                                                        //                .valid
		.cp_data                 (agent_pipeline_008_source0_data),                                                         //                .data
		.cp_startofpacket        (agent_pipeline_008_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (agent_pipeline_008_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (agent_pipeline_008_source0_channel),                                                      //                .channel
		.rf_sink_ready           (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                   //     (terminated)
		.m0_writeresponserequest (),                                                                                        //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                     //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (115),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_startofpacket  (1'b0),                                                                              // (terminated)
		.in_endofpacket    (1'b0),                                                                              // (terminated)
		.out_startofpacket (),                                                                                  // (terminated)
		.out_endofpacket   (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (92),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (103),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (107),
		.PKT_PROTECTION_L          (105),
		.PKT_RESPONSE_STATUS_H     (113),
		.PKT_RESPONSE_STATUS_L     (112),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.ST_CHANNEL_W              (25),
		.ST_DATA_W                 (114),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) audio_fifo_used_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                          //       clk_reset.reset
		.m0_address              (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_010_source0_ready),                                                        //              cp.ready
		.cp_valid                (agent_pipeline_010_source0_valid),                                                        //                .valid
		.cp_data                 (agent_pipeline_010_source0_data),                                                         //                .data
		.cp_startofpacket        (agent_pipeline_010_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (agent_pipeline_010_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (agent_pipeline_010_source0_channel),                                                      //                .channel
		.rf_sink_ready           (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                   //     (terminated)
		.m0_writeresponserequest (),                                                                                        //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                     //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (115),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_startofpacket  (1'b0),                                                                              // (terminated)
		.in_endofpacket    (1'b0),                                                                              // (terminated)
		.out_startofpacket (),                                                                                  // (terminated)
		.out_endofpacket   (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (92),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (103),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (107),
		.PKT_PROTECTION_L          (105),
		.PKT_RESPONSE_STATUS_H     (113),
		.PKT_RESPONSE_STATUS_L     (112),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.ST_CHANNEL_W              (25),
		.ST_DATA_W                 (114),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                    //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_012_source0_ready),                                                           //              cp.ready
		.cp_valid                (agent_pipeline_012_source0_valid),                                                           //                .valid
		.cp_data                 (agent_pipeline_012_source0_data),                                                            //                .data
		.cp_startofpacket        (agent_pipeline_012_source0_startofpacket),                                                   //                .startofpacket
		.cp_endofpacket          (agent_pipeline_012_source0_endofpacket),                                                     //                .endofpacket
		.cp_channel              (agent_pipeline_012_source0_channel),                                                         //                .channel
		.rf_sink_ready           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                      //     (terminated)
		.m0_writeresponserequest (),                                                                                           //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                        //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (115),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                              //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                   // clk_reset.reset
		.in_data           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                 // (terminated)
		.csr_readdata      (),                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                 // (terminated)
		.almost_full_data  (),                                                                                     // (terminated)
		.almost_empty_data (),                                                                                     // (terminated)
		.in_startofpacket  (1'b0),                                                                                 // (terminated)
		.in_endofpacket    (1'b0),                                                                                 // (terminated)
		.out_startofpacket (),                                                                                     // (terminated)
		.out_endofpacket   (),                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                 // (terminated)
		.out_empty         (),                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                 // (terminated)
		.out_error         (),                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                 // (terminated)
		.out_channel       ()                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (92),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (103),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (107),
		.PKT_PROTECTION_L          (105),
		.PKT_RESPONSE_STATUS_H     (113),
		.PKT_RESPONSE_STATUS_L     (112),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.ST_CHANNEL_W              (25),
		.ST_DATA_W                 (114),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                               //       clk_reset.reset
		.m0_address              (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_014_source0_ready),                                                             //              cp.ready
		.cp_valid                (agent_pipeline_014_source0_valid),                                                             //                .valid
		.cp_data                 (agent_pipeline_014_source0_data),                                                              //                .data
		.cp_startofpacket        (agent_pipeline_014_source0_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (agent_pipeline_014_source0_endofpacket),                                                       //                .endofpacket
		.cp_channel              (agent_pipeline_014_source0_channel),                                                           //                .channel
		.rf_sink_ready           (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (115),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                               // clk_reset.reset
		.in_data           (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_startofpacket  (1'b0),                                                                                   // (terminated)
		.in_endofpacket    (1'b0),                                                                                   // (terminated)
		.out_startofpacket (),                                                                                       // (terminated)
		.out_endofpacket   (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (92),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (103),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (107),
		.PKT_PROTECTION_L          (105),
		.PKT_RESPONSE_STATUS_H     (113),
		.PKT_RESPONSE_STATUS_L     (112),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.ST_CHANNEL_W              (25),
		.ST_DATA_W                 (114),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) audio_out_pause_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                          //       clk_reset.reset
		.m0_address              (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_016_source0_ready),                                                        //              cp.ready
		.cp_valid                (agent_pipeline_016_source0_valid),                                                        //                .valid
		.cp_data                 (agent_pipeline_016_source0_data),                                                         //                .data
		.cp_startofpacket        (agent_pipeline_016_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (agent_pipeline_016_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (agent_pipeline_016_source0_channel),                                                      //                .channel
		.rf_sink_ready           (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                   //     (terminated)
		.m0_writeresponserequest (),                                                                                        //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                     //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (115),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_startofpacket  (1'b0),                                                                              // (terminated)
		.in_endofpacket    (1'b0),                                                                              // (terminated)
		.out_startofpacket (),                                                                                  // (terminated)
		.out_endofpacket   (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (92),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (103),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (107),
		.PKT_PROTECTION_L          (105),
		.PKT_RESPONSE_STATUS_H     (113),
		.PKT_RESPONSE_STATUS_L     (112),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.ST_CHANNEL_W              (25),
		.ST_DATA_W                 (114),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) audio_out_stop_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_018_source0_ready),                                                       //              cp.ready
		.cp_valid                (agent_pipeline_018_source0_valid),                                                       //                .valid
		.cp_data                 (agent_pipeline_018_source0_data),                                                        //                .data
		.cp_startofpacket        (agent_pipeline_018_source0_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (agent_pipeline_018_source0_endofpacket),                                                 //                .endofpacket
		.cp_channel              (agent_pipeline_018_source0_channel),                                                     //                .channel
		.rf_sink_ready           (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                  //     (terminated)
		.m0_writeresponserequest (),                                                                                       //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                    //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (115),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.in_data           (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_startofpacket  (1'b0),                                                                             // (terminated)
		.in_endofpacket    (1'b0),                                                                             // (terminated)
		.out_startofpacket (),                                                                                 // (terminated)
		.out_endofpacket   (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (92),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (103),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (107),
		.PKT_PROTECTION_L          (105),
		.PKT_RESPONSE_STATUS_H     (113),
		.PKT_RESPONSE_STATUS_L     (112),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.ST_CHANNEL_W              (25),
		.ST_DATA_W                 (114),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) timer_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                       //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (timer_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_020_source0_ready),                                              //              cp.ready
		.cp_valid                (agent_pipeline_020_source0_valid),                                              //                .valid
		.cp_data                 (agent_pipeline_020_source0_data),                                               //                .data
		.cp_startofpacket        (agent_pipeline_020_source0_startofpacket),                                      //                .startofpacket
		.cp_endofpacket          (agent_pipeline_020_source0_endofpacket),                                        //                .endofpacket
		.cp_channel              (agent_pipeline_020_source0_channel),                                            //                .channel
		.rf_sink_ready           (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (115),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.in_data           (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                          // clk_reset.reset
		.in_data           (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                   // (terminated)
		.csr_read          (1'b0),                                                                    // (terminated)
		.csr_write         (1'b0),                                                                    // (terminated)
		.csr_readdata      (),                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                    // (terminated)
		.almost_full_data  (),                                                                        // (terminated)
		.almost_empty_data (),                                                                        // (terminated)
		.in_startofpacket  (1'b0),                                                                    // (terminated)
		.in_endofpacket    (1'b0),                                                                    // (terminated)
		.out_startofpacket (),                                                                        // (terminated)
		.out_endofpacket   (),                                                                        // (terminated)
		.in_empty          (1'b0),                                                                    // (terminated)
		.out_empty         (),                                                                        // (terminated)
		.in_error          (1'b0),                                                                    // (terminated)
		.out_error         (),                                                                        // (terminated)
		.in_channel        (1'b0),                                                                    // (terminated)
		.out_channel       ()                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (92),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (103),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (107),
		.PKT_PROTECTION_L          (105),
		.PKT_RESPONSE_STATUS_H     (113),
		.PKT_RESPONSE_STATUS_L     (112),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.ST_CHANNEL_W              (25),
		.ST_DATA_W                 (114),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) key_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                     //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (key_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (key_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (key_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (key_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (key_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (key_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (key_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (key_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (key_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (key_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (key_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (key_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (key_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (key_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (key_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (key_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_022_source0_ready),                                            //              cp.ready
		.cp_valid                (agent_pipeline_022_source0_valid),                                            //                .valid
		.cp_data                 (agent_pipeline_022_source0_data),                                             //                .data
		.cp_startofpacket        (agent_pipeline_022_source0_startofpacket),                                    //                .startofpacket
		.cp_endofpacket          (agent_pipeline_022_source0_endofpacket),                                      //                .endofpacket
		.cp_channel              (agent_pipeline_022_source0_channel),                                          //                .channel
		.rf_sink_ready           (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (key_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (key_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (key_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (key_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (key_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (115),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.in_data           (key_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (key_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (key_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (key_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (key_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                       // (terminated)
		.csr_read          (1'b0),                                                                        // (terminated)
		.csr_write         (1'b0),                                                                        // (terminated)
		.csr_readdata      (),                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                        // (terminated)
		.almost_full_data  (),                                                                            // (terminated)
		.almost_empty_data (),                                                                            // (terminated)
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_channel        (1'b0),                                                                        // (terminated)
		.out_channel       ()                                                                             // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.in_data           (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                 // (terminated)
		.csr_read          (1'b0),                                                                  // (terminated)
		.csr_write         (1'b0),                                                                  // (terminated)
		.csr_readdata      (),                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                  // (terminated)
		.almost_full_data  (),                                                                      // (terminated)
		.almost_empty_data (),                                                                      // (terminated)
		.in_startofpacket  (1'b0),                                                                  // (terminated)
		.in_endofpacket    (1'b0),                                                                  // (terminated)
		.out_startofpacket (),                                                                      // (terminated)
		.out_endofpacket   (),                                                                      // (terminated)
		.in_empty          (1'b0),                                                                  // (terminated)
		.out_empty         (),                                                                      // (terminated)
		.in_error          (1'b0),                                                                  // (terminated)
		.out_error         (),                                                                      // (terminated)
		.in_channel        (1'b0),                                                                  // (terminated)
		.out_channel       ()                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (92),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (103),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (107),
		.PKT_PROTECTION_L          (105),
		.PKT_RESPONSE_STATUS_H     (113),
		.PKT_RESPONSE_STATUS_L     (112),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.ST_CHANNEL_W              (25),
		.ST_DATA_W                 (114),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) signal_selector_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                          //       clk_reset.reset
		.m0_address              (signal_selector_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (signal_selector_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (signal_selector_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (signal_selector_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (signal_selector_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (signal_selector_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (signal_selector_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (signal_selector_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (signal_selector_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (signal_selector_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (signal_selector_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (signal_selector_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (signal_selector_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (signal_selector_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (signal_selector_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (signal_selector_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_024_source0_ready),                                                        //              cp.ready
		.cp_valid                (agent_pipeline_024_source0_valid),                                                        //                .valid
		.cp_data                 (agent_pipeline_024_source0_data),                                                         //                .data
		.cp_startofpacket        (agent_pipeline_024_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (agent_pipeline_024_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (agent_pipeline_024_source0_channel),                                                      //                .channel
		.rf_sink_ready           (signal_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (signal_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (signal_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (signal_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (signal_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (signal_selector_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (signal_selector_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (signal_selector_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (signal_selector_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (signal_selector_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (signal_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (signal_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (signal_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (signal_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (signal_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (signal_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                   //     (terminated)
		.m0_writeresponserequest (),                                                                                        //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                     //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (115),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) signal_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (signal_selector_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (signal_selector_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (signal_selector_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (signal_selector_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (signal_selector_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (signal_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (signal_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (signal_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (signal_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (signal_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) signal_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (signal_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (signal_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (signal_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (signal_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (signal_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (signal_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_startofpacket  (1'b0),                                                                              // (terminated)
		.in_endofpacket    (1'b0),                                                                              // (terminated)
		.out_startofpacket (),                                                                                  // (terminated)
		.out_endofpacket   (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (92),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (103),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (107),
		.PKT_PROTECTION_L          (105),
		.PKT_RESPONSE_STATUS_H     (113),
		.PKT_RESPONSE_STATUS_L     (112),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.ST_CHANNEL_W              (25),
		.ST_DATA_W                 (114),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) modulation_selector_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                     //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                              //       clk_reset.reset
		.m0_address              (modulation_selector_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (modulation_selector_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (modulation_selector_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (modulation_selector_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (modulation_selector_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (modulation_selector_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (modulation_selector_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (modulation_selector_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (modulation_selector_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (modulation_selector_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (modulation_selector_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_026_source0_ready),                                                            //              cp.ready
		.cp_valid                (agent_pipeline_026_source0_valid),                                                            //                .valid
		.cp_data                 (agent_pipeline_026_source0_data),                                                             //                .data
		.cp_startofpacket        (agent_pipeline_026_source0_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (agent_pipeline_026_source0_endofpacket),                                                      //                .endofpacket
		.cp_channel              (agent_pipeline_026_source0_channel),                                                          //                .channel
		.rf_sink_ready           (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (115),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) modulation_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.in_data           (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) modulation_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_startofpacket  (1'b0),                                                                                  // (terminated)
		.in_endofpacket    (1'b0),                                                                                  // (terminated)
		.out_startofpacket (),                                                                                      // (terminated)
		.out_endofpacket   (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (92),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (103),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (107),
		.PKT_PROTECTION_L          (105),
		.PKT_RESPONSE_STATUS_H     (113),
		.PKT_RESPONSE_STATUS_L     (112),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.ST_CHANNEL_W              (25),
		.ST_DATA_W                 (114),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) keyboard_keys_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_25_in_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_028_source0_ready),                                                      //              cp.ready
		.cp_valid                (agent_pipeline_028_source0_valid),                                                      //                .valid
		.cp_data                 (agent_pipeline_028_source0_data),                                                       //                .data
		.cp_startofpacket        (agent_pipeline_028_source0_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (agent_pipeline_028_source0_endofpacket),                                                //                .endofpacket
		.cp_channel              (agent_pipeline_028_source0_channel),                                                    //                .channel
		.rf_sink_ready           (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                 //     (terminated)
		.m0_writeresponserequest (),                                                                                      //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                   //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (115),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_25_in_clk),                                                                         //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_25_in_clk),                                                                   //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                              // clk_reset.reset
		.in_data           (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_startofpacket  (1'b0),                                                                            // (terminated)
		.in_endofpacket    (1'b0),                                                                            // (terminated)
		.out_startofpacket (),                                                                                // (terminated)
		.out_endofpacket   (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (92),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (103),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (107),
		.PKT_PROTECTION_L          (105),
		.PKT_RESPONSE_STATUS_H     (113),
		.PKT_RESPONSE_STATUS_L     (112),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.ST_CHANNEL_W              (25),
		.ST_DATA_W                 (114),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) mouse_pos_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_40_in_clk),                                                                     //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (mouse_pos_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (mouse_pos_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (mouse_pos_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (mouse_pos_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (mouse_pos_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (mouse_pos_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (mouse_pos_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (mouse_pos_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (mouse_pos_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (mouse_pos_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (mouse_pos_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_030_source0_ready),                                                  //              cp.ready
		.cp_valid                (agent_pipeline_030_source0_valid),                                                  //                .valid
		.cp_data                 (agent_pipeline_030_source0_data),                                                   //                .data
		.cp_startofpacket        (agent_pipeline_030_source0_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (agent_pipeline_030_source0_endofpacket),                                            //                .endofpacket
		.cp_channel              (agent_pipeline_030_source0_channel),                                                //                .channel
		.rf_sink_ready           (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (115),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) mouse_pos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_40_in_clk),                                                                     //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                // clk_reset.reset
		.in_data           (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) mouse_pos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_40_in_clk),                                                               //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                          // clk_reset.reset
		.in_data           (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                       // (terminated)
		.csr_read          (1'b0),                                                                        // (terminated)
		.csr_write         (1'b0),                                                                        // (terminated)
		.csr_readdata      (),                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                        // (terminated)
		.almost_full_data  (),                                                                            // (terminated)
		.almost_empty_data (),                                                                            // (terminated)
		.in_startofpacket  (1'b0),                                                                        // (terminated)
		.in_endofpacket    (1'b0),                                                                        // (terminated)
		.out_startofpacket (),                                                                            // (terminated)
		.out_endofpacket   (),                                                                            // (terminated)
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_channel        (1'b0),                                                                        // (terminated)
		.out_channel       ()                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (92),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (103),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (107),
		.PKT_PROTECTION_L          (105),
		.PKT_RESPONSE_STATUS_H     (113),
		.PKT_RESPONSE_STATUS_L     (112),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.ST_CHANNEL_W              (25),
		.ST_DATA_W                 (114),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) div_freq_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                   //       clk_reset.reset
		.m0_address              (div_freq_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (div_freq_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (div_freq_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (div_freq_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (div_freq_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (div_freq_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (div_freq_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (div_freq_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (div_freq_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (div_freq_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (div_freq_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (div_freq_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (div_freq_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (div_freq_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (div_freq_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (div_freq_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_032_source0_ready),                                                 //              cp.ready
		.cp_valid                (agent_pipeline_032_source0_valid),                                                 //                .valid
		.cp_data                 (agent_pipeline_032_source0_data),                                                  //                .data
		.cp_startofpacket        (agent_pipeline_032_source0_startofpacket),                                         //                .startofpacket
		.cp_endofpacket          (agent_pipeline_032_source0_endofpacket),                                           //                .endofpacket
		.cp_channel              (agent_pipeline_032_source0_channel),                                               //                .channel
		.rf_sink_ready           (div_freq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (div_freq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (div_freq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (div_freq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (div_freq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (div_freq_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (div_freq_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (div_freq_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (div_freq_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (div_freq_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (div_freq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (div_freq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (div_freq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (div_freq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (div_freq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (div_freq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (115),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) div_freq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.in_data           (div_freq_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (div_freq_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (div_freq_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (div_freq_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (div_freq_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (div_freq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (div_freq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (div_freq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (div_freq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (div_freq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) div_freq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                             // clk_reset.reset
		.in_data           (div_freq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (div_freq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (div_freq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (div_freq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (div_freq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (div_freq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                      // (terminated)
		.csr_read          (1'b0),                                                                       // (terminated)
		.csr_write         (1'b0),                                                                       // (terminated)
		.csr_readdata      (),                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                       // (terminated)
		.almost_full_data  (),                                                                           // (terminated)
		.almost_empty_data (),                                                                           // (terminated)
		.in_startofpacket  (1'b0),                                                                       // (terminated)
		.in_endofpacket    (1'b0),                                                                       // (terminated)
		.out_startofpacket (),                                                                           // (terminated)
		.out_endofpacket   (),                                                                           // (terminated)
		.in_empty          (1'b0),                                                                       // (terminated)
		.out_empty         (),                                                                           // (terminated)
		.in_error          (1'b0),                                                                       // (terminated)
		.out_error         (),                                                                           // (terminated)
		.in_channel        (1'b0),                                                                       // (terminated)
		.out_channel       ()                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (92),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (103),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (107),
		.PKT_PROTECTION_L          (105),
		.PKT_RESPONSE_STATUS_H     (113),
		.PKT_RESPONSE_STATUS_L     (112),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.ST_CHANNEL_W              (25),
		.ST_DATA_W                 (114),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) audio_sel_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (audio_sel_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (audio_sel_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (audio_sel_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (audio_sel_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (audio_sel_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (audio_sel_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (audio_sel_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (audio_sel_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (audio_sel_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (audio_sel_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (audio_sel_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (audio_sel_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (audio_sel_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (audio_sel_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (audio_sel_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (audio_sel_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_034_source0_ready),                                                  //              cp.ready
		.cp_valid                (agent_pipeline_034_source0_valid),                                                  //                .valid
		.cp_data                 (agent_pipeline_034_source0_data),                                                   //                .data
		.cp_startofpacket        (agent_pipeline_034_source0_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (agent_pipeline_034_source0_endofpacket),                                            //                .endofpacket
		.cp_channel              (agent_pipeline_034_source0_channel),                                                //                .channel
		.rf_sink_ready           (audio_sel_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (audio_sel_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (audio_sel_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (audio_sel_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (audio_sel_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (audio_sel_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (audio_sel_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (audio_sel_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (audio_sel_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (audio_sel_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (audio_sel_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (audio_sel_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (audio_sel_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (audio_sel_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (audio_sel_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (audio_sel_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (115),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_sel_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (audio_sel_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (audio_sel_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (audio_sel_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (audio_sel_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (audio_sel_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (audio_sel_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (audio_sel_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (audio_sel_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (audio_sel_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (audio_sel_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_sel_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.in_data           (audio_sel_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (audio_sel_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (audio_sel_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (audio_sel_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (audio_sel_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (audio_sel_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                       // (terminated)
		.csr_read          (1'b0),                                                                        // (terminated)
		.csr_write         (1'b0),                                                                        // (terminated)
		.csr_readdata      (),                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                        // (terminated)
		.almost_full_data  (),                                                                            // (terminated)
		.almost_empty_data (),                                                                            // (terminated)
		.in_startofpacket  (1'b0),                                                                        // (terminated)
		.in_endofpacket    (1'b0),                                                                        // (terminated)
		.out_startofpacket (),                                                                            // (terminated)
		.out_endofpacket   (),                                                                            // (terminated)
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_channel        (1'b0),                                                                        // (terminated)
		.out_channel       ()                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (92),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (103),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (107),
		.PKT_PROTECTION_L          (105),
		.PKT_RESPONSE_STATUS_H     (113),
		.PKT_RESPONSE_STATUS_L     (112),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.ST_CHANNEL_W              (25),
		.ST_DATA_W                 (114),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent (
		.clk                     (cpu_clk_for_sdram_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                                            //       clk_reset.reset
		.m0_address              (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_036_source0_ready),                                                              //              cp.ready
		.cp_valid                (agent_pipeline_036_source0_valid),                                                              //                .valid
		.cp_data                 (agent_pipeline_036_source0_data),                                                               //                .data
		.cp_startofpacket        (agent_pipeline_036_source0_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (agent_pipeline_036_source0_endofpacket),                                                        //                .endofpacket
		.cp_channel              (agent_pipeline_036_source0_channel),                                                            //                .channel
		.rf_sink_ready           (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (115),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (cpu_clk_for_sdram_clk),                                                                         //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                            // clk_reset.reset
		.in_data           (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                          // (terminated)
		.csr_readdata      (),                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                          // (terminated)
		.almost_full_data  (),                                                                                              // (terminated)
		.almost_empty_data (),                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                          // (terminated)
		.out_empty         (),                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                          // (terminated)
		.out_error         (),                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                          // (terminated)
		.out_channel       ()                                                                                               // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (cpu_clk_for_sdram_clk),                                                                   //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                      // clk_reset.reset
		.in_data           (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_startofpacket  (1'b0),                                                                                    // (terminated)
		.in_endofpacket    (1'b0),                                                                                    // (terminated)
		.out_startofpacket (),                                                                                        // (terminated)
		.out_endofpacket   (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (92),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (103),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (107),
		.PKT_PROTECTION_L          (105),
		.PKT_RESPONSE_STATUS_H     (113),
		.PKT_RESPONSE_STATUS_L     (112),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.ST_CHANNEL_W              (25),
		.ST_DATA_W                 (114),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) audio_wrclk_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                             //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                      //       clk_reset.reset
		.m0_address              (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_038_source0_ready),                                                    //              cp.ready
		.cp_valid                (agent_pipeline_038_source0_valid),                                                    //                .valid
		.cp_data                 (agent_pipeline_038_source0_data),                                                     //                .data
		.cp_startofpacket        (agent_pipeline_038_source0_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (agent_pipeline_038_source0_endofpacket),                                              //                .endofpacket
		.cp_channel              (agent_pipeline_038_source0_channel),                                                  //                .channel
		.rf_sink_ready           (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (115),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                      // clk_reset.reset
		.in_data           (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.in_data           (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_startofpacket  (1'b0),                                                                          // (terminated)
		.in_endofpacket    (1'b0),                                                                          // (terminated)
		.out_startofpacket (),                                                                              // (terminated)
		.out_endofpacket   (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (92),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (103),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (107),
		.PKT_PROTECTION_L          (105),
		.PKT_RESPONSE_STATUS_H     (113),
		.PKT_RESPONSE_STATUS_L     (112),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.ST_CHANNEL_W              (25),
		.ST_DATA_W                 (114),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) audio_wrreq_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                             //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                      //       clk_reset.reset
		.m0_address              (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_040_source0_ready),                                                    //              cp.ready
		.cp_valid                (agent_pipeline_040_source0_valid),                                                    //                .valid
		.cp_data                 (agent_pipeline_040_source0_data),                                                     //                .data
		.cp_startofpacket        (agent_pipeline_040_source0_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (agent_pipeline_040_source0_endofpacket),                                              //                .endofpacket
		.cp_channel              (agent_pipeline_040_source0_channel),                                                  //                .channel
		.rf_sink_ready           (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (115),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                      // clk_reset.reset
		.in_data           (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.in_data           (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_startofpacket  (1'b0),                                                                          // (terminated)
		.in_endofpacket    (1'b0),                                                                          // (terminated)
		.out_startofpacket (),                                                                              // (terminated)
		.out_endofpacket   (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (74),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (80),
		.PKT_SRC_ID_L              (76),
		.PKT_DEST_ID_H             (85),
		.PKT_DEST_ID_L             (81),
		.PKT_BURSTWRAP_H           (66),
		.PKT_BURSTWRAP_L           (64),
		.PKT_BYTE_CNT_H            (63),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (89),
		.PKT_PROTECTION_L          (87),
		.PKT_RESPONSE_STATUS_H     (95),
		.PKT_RESPONSE_STATUS_L     (94),
		.PKT_BURST_SIZE_H          (69),
		.PKT_BURST_SIZE_L          (67),
		.ST_CHANNEL_W              (25),
		.ST_DATA_W                 (96),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (cpu_clk_for_sdram_clk),                                                         //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                            //       clk_reset.reset
		.m0_address              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_042_source0_ready),                                              //              cp.ready
		.cp_valid                (agent_pipeline_042_source0_valid),                                              //                .valid
		.cp_data                 (agent_pipeline_042_source0_data),                                               //                .data
		.cp_startofpacket        (agent_pipeline_042_source0_startofpacket),                                      //                .startofpacket
		.cp_endofpacket          (agent_pipeline_042_source0_endofpacket),                                        //                .endofpacket
		.cp_channel              (agent_pipeline_042_source0_channel),                                            //                .channel
		.rf_sink_ready           (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (97),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (cpu_clk_for_sdram_clk),                                                         //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                            // clk_reset.reset
		.in_data           (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (18),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (cpu_clk_for_sdram_clk),                                                   //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                      // clk_reset.reset
		.in_data           (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                   // (terminated)
		.csr_read          (1'b0),                                                                    // (terminated)
		.csr_write         (1'b0),                                                                    // (terminated)
		.csr_readdata      (),                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                    // (terminated)
		.almost_full_data  (),                                                                        // (terminated)
		.almost_empty_data (),                                                                        // (terminated)
		.in_startofpacket  (1'b0),                                                                    // (terminated)
		.in_endofpacket    (1'b0),                                                                    // (terminated)
		.out_startofpacket (),                                                                        // (terminated)
		.out_endofpacket   (),                                                                        // (terminated)
		.in_empty          (1'b0),                                                                    // (terminated)
		.out_empty         (),                                                                        // (terminated)
		.in_error          (1'b0),                                                                    // (terminated)
		.out_error         (),                                                                        // (terminated)
		.in_channel        (1'b0),                                                                    // (terminated)
		.out_channel       ()                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (92),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (103),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (107),
		.PKT_PROTECTION_L          (105),
		.PKT_RESPONSE_STATUS_H     (113),
		.PKT_RESPONSE_STATUS_L     (112),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.ST_CHANNEL_W              (25),
		.ST_DATA_W                 (114),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                 //       clk_reset.reset
		.m0_address              (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_044_source0_ready),                                                               //              cp.ready
		.cp_valid                (agent_pipeline_044_source0_valid),                                                               //                .valid
		.cp_data                 (agent_pipeline_044_source0_data),                                                                //                .data
		.cp_startofpacket        (agent_pipeline_044_source0_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (agent_pipeline_044_source0_endofpacket),                                                         //                .endofpacket
		.cp_channel              (agent_pipeline_044_source0_channel),                                                             //                .channel
		.rf_sink_ready           (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (115),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                 // clk_reset.reset
		.in_data           (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                          // (terminated)
		.csr_read          (1'b0),                                                                                           // (terminated)
		.csr_write         (1'b0),                                                                                           // (terminated)
		.csr_readdata      (),                                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                           // (terminated)
		.almost_full_data  (),                                                                                               // (terminated)
		.almost_empty_data (),                                                                                               // (terminated)
		.in_empty          (1'b0),                                                                                           // (terminated)
		.out_empty         (),                                                                                               // (terminated)
		.in_error          (1'b0),                                                                                           // (terminated)
		.out_error         (),                                                                                               // (terminated)
		.in_channel        (1'b0),                                                                                           // (terminated)
		.out_channel       ()                                                                                                // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_startofpacket  (1'b0),                                                                                     // (terminated)
		.in_endofpacket    (1'b0),                                                                                     // (terminated)
		.out_startofpacket (),                                                                                         // (terminated)
		.out_endofpacket   (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (92),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (103),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (107),
		.PKT_PROTECTION_L          (105),
		.PKT_RESPONSE_STATUS_H     (113),
		.PKT_RESPONSE_STATUS_L     (112),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.ST_CHANNEL_W              (25),
		.ST_DATA_W                 (114),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) lfsr_val_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                   //       clk_reset.reset
		.m0_address              (lfsr_val_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (lfsr_val_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (lfsr_val_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (lfsr_val_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (lfsr_val_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (lfsr_val_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (lfsr_val_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (lfsr_val_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (lfsr_val_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (lfsr_val_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (lfsr_val_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_046_source0_ready),                                                 //              cp.ready
		.cp_valid                (agent_pipeline_046_source0_valid),                                                 //                .valid
		.cp_data                 (agent_pipeline_046_source0_data),                                                  //                .data
		.cp_startofpacket        (agent_pipeline_046_source0_startofpacket),                                         //                .startofpacket
		.cp_endofpacket          (agent_pipeline_046_source0_endofpacket),                                           //                .endofpacket
		.cp_channel              (agent_pipeline_046_source0_channel),                                               //                .channel
		.rf_sink_ready           (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (115),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) lfsr_val_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.in_data           (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) lfsr_val_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                             // clk_reset.reset
		.in_data           (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                      // (terminated)
		.csr_read          (1'b0),                                                                       // (terminated)
		.csr_write         (1'b0),                                                                       // (terminated)
		.csr_readdata      (),                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                       // (terminated)
		.almost_full_data  (),                                                                           // (terminated)
		.almost_empty_data (),                                                                           // (terminated)
		.in_startofpacket  (1'b0),                                                                       // (terminated)
		.in_endofpacket    (1'b0),                                                                       // (terminated)
		.out_startofpacket (),                                                                           // (terminated)
		.out_endofpacket   (),                                                                           // (terminated)
		.in_empty          (1'b0),                                                                       // (terminated)
		.out_empty         (),                                                                           // (terminated)
		.in_error          (1'b0),                                                                       // (terminated)
		.out_error         (),                                                                           // (terminated)
		.in_channel        (1'b0),                                                                       // (terminated)
		.out_channel       ()                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (92),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (98),
		.PKT_SRC_ID_L              (94),
		.PKT_DEST_ID_H             (103),
		.PKT_DEST_ID_L             (99),
		.PKT_BURSTWRAP_H           (84),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (107),
		.PKT_PROTECTION_L          (105),
		.PKT_RESPONSE_STATUS_H     (113),
		.PKT_RESPONSE_STATUS_L     (112),
		.PKT_BURST_SIZE_H          (87),
		.PKT_BURST_SIZE_L          (85),
		.ST_CHANNEL_W              (25),
		.ST_DATA_W                 (114),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) dds_increment_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (dds_increment_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (dds_increment_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (dds_increment_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (dds_increment_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (dds_increment_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (dds_increment_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (dds_increment_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (dds_increment_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (dds_increment_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (dds_increment_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (dds_increment_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (dds_increment_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (dds_increment_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (dds_increment_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (dds_increment_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (dds_increment_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (agent_pipeline_048_source0_ready),                                                      //              cp.ready
		.cp_valid                (agent_pipeline_048_source0_valid),                                                      //                .valid
		.cp_data                 (agent_pipeline_048_source0_data),                                                       //                .data
		.cp_startofpacket        (agent_pipeline_048_source0_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (agent_pipeline_048_source0_endofpacket),                                                //                .endofpacket
		.cp_channel              (agent_pipeline_048_source0_channel),                                                    //                .channel
		.rf_sink_ready           (dds_increment_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (dds_increment_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (dds_increment_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (dds_increment_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (dds_increment_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (dds_increment_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (dds_increment_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (dds_increment_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (dds_increment_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (dds_increment_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (dds_increment_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (dds_increment_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (dds_increment_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (dds_increment_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (dds_increment_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (dds_increment_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                 //     (terminated)
		.m0_writeresponserequest (),                                                                                      //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                   //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (115),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dds_increment_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (dds_increment_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (dds_increment_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (dds_increment_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (dds_increment_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (dds_increment_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (dds_increment_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (dds_increment_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (dds_increment_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (dds_increment_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (dds_increment_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dds_increment_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (dds_increment_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (dds_increment_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (dds_increment_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (dds_increment_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (dds_increment_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (dds_increment_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_startofpacket  (1'b0),                                                                            // (terminated)
		.in_endofpacket    (1'b0),                                                                            // (terminated)
		.out_startofpacket (),                                                                                // (terminated)
		.out_endofpacket   (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	DE2_QSYS_addr_router addr_router (
		.sink_ready         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                     //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                       //       src.ready
		.src_valid          (addr_router_src_valid),                                                       //          .valid
		.src_data           (addr_router_src_data),                                                        //          .data
		.src_channel        (addr_router_src_channel),                                                     //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                  //          .endofpacket
	);

	DE2_QSYS_addr_router_001 addr_router_001 (
		.sink_ready         (vga_to_sdram_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (vga_to_sdram_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (vga_to_sdram_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (vga_to_sdram_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (vga_to_sdram_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (cpu_clk_for_sdram_clk),                                                    //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                //          .valid
		.src_data           (addr_router_001_src_data),                                                 //          .data
		.src_channel        (addr_router_001_src_channel),                                              //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                           //          .endofpacket
	);

	DE2_QSYS_addr_router_002 addr_router_002 (
		.sink_ready         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                          //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                          //          .valid
		.src_data           (addr_router_002_src_data),                                                           //          .data
		.src_channel        (addr_router_002_src_channel),                                                        //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                                  //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                                     //          .endofpacket
	);

	DE2_QSYS_id_router id_router (
		.sink_ready         (agent_pipeline_001_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_001_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_001_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_001_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_001_source0_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),           // clk_reset.reset
		.src_ready          (id_router_src_ready),                      //       src.ready
		.src_valid          (id_router_src_valid),                      //          .valid
		.src_data           (id_router_src_data),                       //          .data
		.src_channel        (id_router_src_channel),                    //          .channel
		.src_startofpacket  (id_router_src_startofpacket),              //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                 //          .endofpacket
	);

	DE2_QSYS_id_router id_router_001 (
		.sink_ready         (agent_pipeline_003_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_003_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_003_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_003_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_003_source0_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),           // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                  //       src.ready
		.src_valid          (id_router_001_src_valid),                  //          .valid
		.src_data           (id_router_001_src_data),                   //          .data
		.src_channel        (id_router_001_src_channel),                //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)             //          .endofpacket
	);

	DE2_QSYS_id_router id_router_002 (
		.sink_ready         (agent_pipeline_005_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_005_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_005_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_005_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_005_source0_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),           // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                  //       src.ready
		.src_valid          (id_router_002_src_valid),                  //          .valid
		.src_data           (id_router_002_src_data),                   //          .data
		.src_channel        (id_router_002_src_channel),                //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)             //          .endofpacket
	);

	DE2_QSYS_id_router id_router_003 (
		.sink_ready         (agent_pipeline_007_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_007_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_007_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_007_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_007_source0_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),           // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                  //       src.ready
		.src_valid          (id_router_003_src_valid),                  //          .valid
		.src_data           (id_router_003_src_data),                   //          .data
		.src_channel        (id_router_003_src_channel),                //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)             //          .endofpacket
	);

	DE2_QSYS_id_router id_router_004 (
		.sink_ready         (agent_pipeline_009_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_009_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_009_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_009_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_009_source0_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),           // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                  //       src.ready
		.src_valid          (id_router_004_src_valid),                  //          .valid
		.src_data           (id_router_004_src_data),                   //          .data
		.src_channel        (id_router_004_src_channel),                //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)             //          .endofpacket
	);

	DE2_QSYS_id_router id_router_005 (
		.sink_ready         (agent_pipeline_011_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_011_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_011_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_011_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_011_source0_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),           // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                  //       src.ready
		.src_valid          (id_router_005_src_valid),                  //          .valid
		.src_data           (id_router_005_src_data),                   //          .data
		.src_channel        (id_router_005_src_channel),                //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)             //          .endofpacket
	);

	DE2_QSYS_id_router_006 id_router_006 (
		.sink_ready         (agent_pipeline_013_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_013_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_013_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_013_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_013_source0_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),       // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                  //       src.ready
		.src_valid          (id_router_006_src_valid),                  //          .valid
		.src_data           (id_router_006_src_data),                   //          .data
		.src_channel        (id_router_006_src_channel),                //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)             //          .endofpacket
	);

	DE2_QSYS_id_router id_router_007 (
		.sink_ready         (agent_pipeline_015_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_015_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_015_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_015_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_015_source0_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),           // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                  //       src.ready
		.src_valid          (id_router_007_src_valid),                  //          .valid
		.src_data           (id_router_007_src_data),                   //          .data
		.src_channel        (id_router_007_src_channel),                //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)             //          .endofpacket
	);

	DE2_QSYS_id_router id_router_008 (
		.sink_ready         (agent_pipeline_017_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_017_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_017_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_017_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_017_source0_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),           // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                  //       src.ready
		.src_valid          (id_router_008_src_valid),                  //          .valid
		.src_data           (id_router_008_src_data),                   //          .data
		.src_channel        (id_router_008_src_channel),                //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)             //          .endofpacket
	);

	DE2_QSYS_id_router id_router_009 (
		.sink_ready         (agent_pipeline_019_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_019_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_019_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_019_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_019_source0_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),           // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                  //       src.ready
		.src_valid          (id_router_009_src_valid),                  //          .valid
		.src_data           (id_router_009_src_data),                   //          .data
		.src_channel        (id_router_009_src_channel),                //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)             //          .endofpacket
	);

	DE2_QSYS_id_router id_router_010 (
		.sink_ready         (agent_pipeline_021_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_021_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_021_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_021_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_021_source0_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),           // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                  //       src.ready
		.src_valid          (id_router_010_src_valid),                  //          .valid
		.src_data           (id_router_010_src_data),                   //          .data
		.src_channel        (id_router_010_src_channel),                //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)             //          .endofpacket
	);

	DE2_QSYS_id_router id_router_011 (
		.sink_ready         (agent_pipeline_023_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_023_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_023_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_023_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_023_source0_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),           // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                  //       src.ready
		.src_valid          (id_router_011_src_valid),                  //          .valid
		.src_data           (id_router_011_src_data),                   //          .data
		.src_channel        (id_router_011_src_channel),                //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)             //          .endofpacket
	);

	DE2_QSYS_id_router id_router_012 (
		.sink_ready         (agent_pipeline_025_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_025_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_025_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_025_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_025_source0_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),           // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                  //       src.ready
		.src_valid          (id_router_012_src_valid),                  //          .valid
		.src_data           (id_router_012_src_data),                   //          .data
		.src_channel        (id_router_012_src_channel),                //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)             //          .endofpacket
	);

	DE2_QSYS_id_router id_router_013 (
		.sink_ready         (agent_pipeline_027_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_027_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_027_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_027_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_027_source0_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),           // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                  //       src.ready
		.src_valid          (id_router_013_src_valid),                  //          .valid
		.src_data           (id_router_013_src_data),                   //          .data
		.src_channel        (id_router_013_src_channel),                //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)             //          .endofpacket
	);

	DE2_QSYS_id_router id_router_014 (
		.sink_ready         (agent_pipeline_029_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_029_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_029_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_029_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_029_source0_endofpacket),   //          .endofpacket
		.clk                (clk_25_in_clk),                            //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),       // clk_reset.reset
		.src_ready          (id_router_014_src_ready),                  //       src.ready
		.src_valid          (id_router_014_src_valid),                  //          .valid
		.src_data           (id_router_014_src_data),                   //          .data
		.src_channel        (id_router_014_src_channel),                //          .channel
		.src_startofpacket  (id_router_014_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_014_src_endofpacket)             //          .endofpacket
	);

	DE2_QSYS_id_router id_router_015 (
		.sink_ready         (agent_pipeline_031_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_031_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_031_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_031_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_031_source0_endofpacket),   //          .endofpacket
		.clk                (clk_40_in_clk),                            //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),       // clk_reset.reset
		.src_ready          (id_router_015_src_ready),                  //       src.ready
		.src_valid          (id_router_015_src_valid),                  //          .valid
		.src_data           (id_router_015_src_data),                   //          .data
		.src_channel        (id_router_015_src_channel),                //          .channel
		.src_startofpacket  (id_router_015_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_015_src_endofpacket)             //          .endofpacket
	);

	DE2_QSYS_id_router id_router_016 (
		.sink_ready         (agent_pipeline_033_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_033_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_033_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_033_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_033_source0_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),           // clk_reset.reset
		.src_ready          (id_router_016_src_ready),                  //       src.ready
		.src_valid          (id_router_016_src_valid),                  //          .valid
		.src_data           (id_router_016_src_data),                   //          .data
		.src_channel        (id_router_016_src_channel),                //          .channel
		.src_startofpacket  (id_router_016_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_016_src_endofpacket)             //          .endofpacket
	);

	DE2_QSYS_id_router id_router_017 (
		.sink_ready         (agent_pipeline_035_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_035_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_035_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_035_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_035_source0_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),           // clk_reset.reset
		.src_ready          (id_router_017_src_ready),                  //       src.ready
		.src_valid          (id_router_017_src_valid),                  //          .valid
		.src_data           (id_router_017_src_data),                   //          .data
		.src_channel        (id_router_017_src_channel),                //          .channel
		.src_startofpacket  (id_router_017_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_017_src_endofpacket)             //          .endofpacket
	);

	DE2_QSYS_id_router id_router_018 (
		.sink_ready         (agent_pipeline_037_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_037_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_037_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_037_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_037_source0_endofpacket),   //          .endofpacket
		.clk                (cpu_clk_for_sdram_clk),                    //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),       // clk_reset.reset
		.src_ready          (id_router_018_src_ready),                  //       src.ready
		.src_valid          (id_router_018_src_valid),                  //          .valid
		.src_data           (id_router_018_src_data),                   //          .data
		.src_channel        (id_router_018_src_channel),                //          .channel
		.src_startofpacket  (id_router_018_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_018_src_endofpacket)             //          .endofpacket
	);

	DE2_QSYS_id_router id_router_019 (
		.sink_ready         (agent_pipeline_039_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_039_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_039_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_039_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_039_source0_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),           // clk_reset.reset
		.src_ready          (id_router_019_src_ready),                  //       src.ready
		.src_valid          (id_router_019_src_valid),                  //          .valid
		.src_data           (id_router_019_src_data),                   //          .data
		.src_channel        (id_router_019_src_channel),                //          .channel
		.src_startofpacket  (id_router_019_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_019_src_endofpacket)             //          .endofpacket
	);

	DE2_QSYS_id_router id_router_020 (
		.sink_ready         (agent_pipeline_041_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_041_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_041_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_041_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_041_source0_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),           // clk_reset.reset
		.src_ready          (id_router_020_src_ready),                  //       src.ready
		.src_valid          (id_router_020_src_valid),                  //          .valid
		.src_data           (id_router_020_src_data),                   //          .data
		.src_channel        (id_router_020_src_channel),                //          .channel
		.src_startofpacket  (id_router_020_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_020_src_endofpacket)             //          .endofpacket
	);

	DE2_QSYS_id_router_021 id_router_021 (
		.sink_ready         (agent_pipeline_043_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_043_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_043_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_043_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_043_source0_endofpacket),   //          .endofpacket
		.clk                (cpu_clk_for_sdram_clk),                    //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),       // clk_reset.reset
		.src_ready          (id_router_021_src_ready),                  //       src.ready
		.src_valid          (id_router_021_src_valid),                  //          .valid
		.src_data           (id_router_021_src_data),                   //          .data
		.src_channel        (id_router_021_src_channel),                //          .channel
		.src_startofpacket  (id_router_021_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_021_src_endofpacket)             //          .endofpacket
	);

	DE2_QSYS_id_router id_router_022 (
		.sink_ready         (agent_pipeline_045_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_045_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_045_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_045_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_045_source0_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),           // clk_reset.reset
		.src_ready          (id_router_022_src_ready),                  //       src.ready
		.src_valid          (id_router_022_src_valid),                  //          .valid
		.src_data           (id_router_022_src_data),                   //          .data
		.src_channel        (id_router_022_src_channel),                //          .channel
		.src_startofpacket  (id_router_022_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_022_src_endofpacket)             //          .endofpacket
	);

	DE2_QSYS_id_router id_router_023 (
		.sink_ready         (agent_pipeline_047_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_047_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_047_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_047_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_047_source0_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),           // clk_reset.reset
		.src_ready          (id_router_023_src_ready),                  //       src.ready
		.src_valid          (id_router_023_src_valid),                  //          .valid
		.src_data           (id_router_023_src_data),                   //          .data
		.src_channel        (id_router_023_src_channel),                //          .channel
		.src_startofpacket  (id_router_023_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_023_src_endofpacket)             //          .endofpacket
	);

	DE2_QSYS_id_router id_router_024 (
		.sink_ready         (agent_pipeline_049_source0_ready),         //      sink.ready
		.sink_valid         (agent_pipeline_049_source0_valid),         //          .valid
		.sink_data          (agent_pipeline_049_source0_data),          //          .data
		.sink_startofpacket (agent_pipeline_049_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (agent_pipeline_049_source0_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),           // clk_reset.reset
		.src_ready          (id_router_024_src_ready),                  //       src.ready
		.src_valid          (id_router_024_src_valid),                  //          .valid
		.src_data           (id_router_024_src_data),                   //          .data
		.src_channel        (id_router_024_src_channel),                //          .channel
		.src_startofpacket  (id_router_024_src_startofpacket),          //          .startofpacket
		.src_endofpacket    (id_router_024_src_endofpacket)             //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (103),
		.PKT_DEST_ID_L             (99),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.MAX_OUTSTANDING_RESPONSES (21),
		.PIPELINED                 (0),
		.ST_DATA_W                 (114),
		.ST_CHANNEL_W              (25),
		.VALID_WIDTH               (1),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (clk_clk),                                    //       clk.clk
		.reset                  (rst_controller_001_reset_out_reset),         // clk_reset.reset
		.cmd_sink_ready         (addr_router_002_src_ready),                  //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_002_src_valid),                  //          .valid
		.cmd_sink_data          (addr_router_002_src_data),                   //          .data
		.cmd_sink_channel       (addr_router_002_src_channel),                //          .channel
		.cmd_sink_startofpacket (addr_router_002_src_startofpacket),          //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_002_src_endofpacket),            //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),                      //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),                       //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),                    //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),              //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),                //          .endofpacket
		.cmd_src_valid          (limiter_cmd_src_valid),                      //          .valid
		.rsp_sink_ready         (limiter_pipeline_001_source0_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (limiter_pipeline_001_source0_valid),         //          .valid
		.rsp_sink_channel       (limiter_pipeline_001_source0_channel),       //          .channel
		.rsp_sink_data          (limiter_pipeline_001_source0_data),          //          .data
		.rsp_sink_startofpacket (limiter_pipeline_001_source0_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (limiter_pipeline_001_source0_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),                      //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),                      //          .valid
		.rsp_src_data           (limiter_rsp_src_data),                       //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),                    //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),              //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket)                 //          .endofpacket
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (74),
		.PKT_BYTE_CNT_H            (63),
		.PKT_BYTE_CNT_L            (56),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (69),
		.PKT_BURST_SIZE_L          (67),
		.PKT_BURST_TYPE_H          (71),
		.PKT_BURST_TYPE_L          (70),
		.PKT_BURSTWRAP_H           (66),
		.PKT_BURSTWRAP_L           (64),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (96),
		.ST_CHANNEL_W              (25),
		.OUT_BYTE_CNT_H            (57),
		.OUT_BURSTWRAP_H           (66),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter (
		.clk                   (cpu_clk_for_sdram_clk),               //       cr0.clk
		.reset                 (rst_controller_004_reset_out_reset),  // cr0_reset.reset
		.sink0_valid           (width_adapter_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_src_data),              //          .data
		.sink0_channel         (width_adapter_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_src_ready),             //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (clk_clk),                        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req  (),                               // (terminated)
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.reset_in1  (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk        (clk_clk),                            //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_002 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (clk_25_in_clk),                      //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_003 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (clk_40_in_clk),                      //       clk.clk
		.reset_out  (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_004 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (cpu_clk_for_sdram_clk),              //       clk.clk
		.reset_out  (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	DE2_QSYS_cmd_xbar_demux cmd_xbar_demux (
		.clk                 (clk_clk),                            //       clk.clk
		.reset               (rst_controller_001_reset_out_reset), // clk_reset.reset
		.sink_ready          (addr_router_src_ready),              //      sink.ready
		.sink_channel        (addr_router_src_channel),            //          .channel
		.sink_data           (addr_router_src_data),               //          .data
		.sink_startofpacket  (addr_router_src_startofpacket),      //          .startofpacket
		.sink_endofpacket    (addr_router_src_endofpacket),        //          .endofpacket
		.sink_valid          (addr_router_src_valid),              //          .valid
		.src0_ready          (cmd_xbar_demux_src0_ready),          //      src0.ready
		.src0_valid          (cmd_xbar_demux_src0_valid),          //          .valid
		.src0_data           (cmd_xbar_demux_src0_data),           //          .data
		.src0_channel        (cmd_xbar_demux_src0_channel),        //          .channel
		.src0_startofpacket  (cmd_xbar_demux_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_src0_endofpacket),    //          .endofpacket
		.src1_ready          (cmd_xbar_demux_src1_ready),          //      src1.ready
		.src1_valid          (cmd_xbar_demux_src1_valid),          //          .valid
		.src1_data           (cmd_xbar_demux_src1_data),           //          .data
		.src1_channel        (cmd_xbar_demux_src1_channel),        //          .channel
		.src1_startofpacket  (cmd_xbar_demux_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_src1_endofpacket),    //          .endofpacket
		.src2_ready          (cmd_xbar_demux_src2_ready),          //      src2.ready
		.src2_valid          (cmd_xbar_demux_src2_valid),          //          .valid
		.src2_data           (cmd_xbar_demux_src2_data),           //          .data
		.src2_channel        (cmd_xbar_demux_src2_channel),        //          .channel
		.src2_startofpacket  (cmd_xbar_demux_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_src2_endofpacket),    //          .endofpacket
		.src3_ready          (cmd_xbar_demux_src3_ready),          //      src3.ready
		.src3_valid          (cmd_xbar_demux_src3_valid),          //          .valid
		.src3_data           (cmd_xbar_demux_src3_data),           //          .data
		.src3_channel        (cmd_xbar_demux_src3_channel),        //          .channel
		.src3_startofpacket  (cmd_xbar_demux_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_src3_endofpacket),    //          .endofpacket
		.src4_ready          (cmd_xbar_demux_src4_ready),          //      src4.ready
		.src4_valid          (cmd_xbar_demux_src4_valid),          //          .valid
		.src4_data           (cmd_xbar_demux_src4_data),           //          .data
		.src4_channel        (cmd_xbar_demux_src4_channel),        //          .channel
		.src4_startofpacket  (cmd_xbar_demux_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_src4_endofpacket),    //          .endofpacket
		.src5_ready          (cmd_xbar_demux_src5_ready),          //      src5.ready
		.src5_valid          (cmd_xbar_demux_src5_valid),          //          .valid
		.src5_data           (cmd_xbar_demux_src5_data),           //          .data
		.src5_channel        (cmd_xbar_demux_src5_channel),        //          .channel
		.src5_startofpacket  (cmd_xbar_demux_src5_startofpacket),  //          .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_src5_endofpacket),    //          .endofpacket
		.src6_ready          (cmd_xbar_demux_src6_ready),          //      src6.ready
		.src6_valid          (cmd_xbar_demux_src6_valid),          //          .valid
		.src6_data           (cmd_xbar_demux_src6_data),           //          .data
		.src6_channel        (cmd_xbar_demux_src6_channel),        //          .channel
		.src6_startofpacket  (cmd_xbar_demux_src6_startofpacket),  //          .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_src6_endofpacket),    //          .endofpacket
		.src7_ready          (cmd_xbar_demux_src7_ready),          //      src7.ready
		.src7_valid          (cmd_xbar_demux_src7_valid),          //          .valid
		.src7_data           (cmd_xbar_demux_src7_data),           //          .data
		.src7_channel        (cmd_xbar_demux_src7_channel),        //          .channel
		.src7_startofpacket  (cmd_xbar_demux_src7_startofpacket),  //          .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_src7_endofpacket),    //          .endofpacket
		.src8_ready          (cmd_xbar_demux_src8_ready),          //      src8.ready
		.src8_valid          (cmd_xbar_demux_src8_valid),          //          .valid
		.src8_data           (cmd_xbar_demux_src8_data),           //          .data
		.src8_channel        (cmd_xbar_demux_src8_channel),        //          .channel
		.src8_startofpacket  (cmd_xbar_demux_src8_startofpacket),  //          .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_src8_endofpacket),    //          .endofpacket
		.src9_ready          (cmd_xbar_demux_src9_ready),          //      src9.ready
		.src9_valid          (cmd_xbar_demux_src9_valid),          //          .valid
		.src9_data           (cmd_xbar_demux_src9_data),           //          .data
		.src9_channel        (cmd_xbar_demux_src9_channel),        //          .channel
		.src9_startofpacket  (cmd_xbar_demux_src9_startofpacket),  //          .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_src9_endofpacket),    //          .endofpacket
		.src10_ready         (cmd_xbar_demux_src10_ready),         //     src10.ready
		.src10_valid         (cmd_xbar_demux_src10_valid),         //          .valid
		.src10_data          (cmd_xbar_demux_src10_data),          //          .data
		.src10_channel       (cmd_xbar_demux_src10_channel),       //          .channel
		.src10_startofpacket (cmd_xbar_demux_src10_startofpacket), //          .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_src10_endofpacket),   //          .endofpacket
		.src11_ready         (cmd_xbar_demux_src11_ready),         //     src11.ready
		.src11_valid         (cmd_xbar_demux_src11_valid),         //          .valid
		.src11_data          (cmd_xbar_demux_src11_data),          //          .data
		.src11_channel       (cmd_xbar_demux_src11_channel),       //          .channel
		.src11_startofpacket (cmd_xbar_demux_src11_startofpacket), //          .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_src11_endofpacket),   //          .endofpacket
		.src12_ready         (cmd_xbar_demux_src12_ready),         //     src12.ready
		.src12_valid         (cmd_xbar_demux_src12_valid),         //          .valid
		.src12_data          (cmd_xbar_demux_src12_data),          //          .data
		.src12_channel       (cmd_xbar_demux_src12_channel),       //          .channel
		.src12_startofpacket (cmd_xbar_demux_src12_startofpacket), //          .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_src12_endofpacket),   //          .endofpacket
		.src13_ready         (cmd_xbar_demux_src13_ready),         //     src13.ready
		.src13_valid         (cmd_xbar_demux_src13_valid),         //          .valid
		.src13_data          (cmd_xbar_demux_src13_data),          //          .data
		.src13_channel       (cmd_xbar_demux_src13_channel),       //          .channel
		.src13_startofpacket (cmd_xbar_demux_src13_startofpacket), //          .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_src13_endofpacket),   //          .endofpacket
		.src14_ready         (cmd_xbar_demux_src14_ready),         //     src14.ready
		.src14_valid         (cmd_xbar_demux_src14_valid),         //          .valid
		.src14_data          (cmd_xbar_demux_src14_data),          //          .data
		.src14_channel       (cmd_xbar_demux_src14_channel),       //          .channel
		.src14_startofpacket (cmd_xbar_demux_src14_startofpacket), //          .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_src14_endofpacket),   //          .endofpacket
		.src15_ready         (cmd_xbar_demux_src15_ready),         //     src15.ready
		.src15_valid         (cmd_xbar_demux_src15_valid),         //          .valid
		.src15_data          (cmd_xbar_demux_src15_data),          //          .data
		.src15_channel       (cmd_xbar_demux_src15_channel),       //          .channel
		.src15_startofpacket (cmd_xbar_demux_src15_startofpacket), //          .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_src15_endofpacket),   //          .endofpacket
		.src16_ready         (cmd_xbar_demux_src16_ready),         //     src16.ready
		.src16_valid         (cmd_xbar_demux_src16_valid),         //          .valid
		.src16_data          (cmd_xbar_demux_src16_data),          //          .data
		.src16_channel       (cmd_xbar_demux_src16_channel),       //          .channel
		.src16_startofpacket (cmd_xbar_demux_src16_startofpacket), //          .startofpacket
		.src16_endofpacket   (cmd_xbar_demux_src16_endofpacket),   //          .endofpacket
		.src17_ready         (cmd_xbar_demux_src17_ready),         //     src17.ready
		.src17_valid         (cmd_xbar_demux_src17_valid),         //          .valid
		.src17_data          (cmd_xbar_demux_src17_data),          //          .data
		.src17_channel       (cmd_xbar_demux_src17_channel),       //          .channel
		.src17_startofpacket (cmd_xbar_demux_src17_startofpacket), //          .startofpacket
		.src17_endofpacket   (cmd_xbar_demux_src17_endofpacket),   //          .endofpacket
		.src18_ready         (cmd_xbar_demux_src18_ready),         //     src18.ready
		.src18_valid         (cmd_xbar_demux_src18_valid),         //          .valid
		.src18_data          (cmd_xbar_demux_src18_data),          //          .data
		.src18_channel       (cmd_xbar_demux_src18_channel),       //          .channel
		.src18_startofpacket (cmd_xbar_demux_src18_startofpacket), //          .startofpacket
		.src18_endofpacket   (cmd_xbar_demux_src18_endofpacket),   //          .endofpacket
		.src19_ready         (cmd_xbar_demux_src19_ready),         //     src19.ready
		.src19_valid         (cmd_xbar_demux_src19_valid),         //          .valid
		.src19_data          (cmd_xbar_demux_src19_data),          //          .data
		.src19_channel       (cmd_xbar_demux_src19_channel),       //          .channel
		.src19_startofpacket (cmd_xbar_demux_src19_startofpacket), //          .startofpacket
		.src19_endofpacket   (cmd_xbar_demux_src19_endofpacket),   //          .endofpacket
		.src20_ready         (cmd_xbar_demux_src20_ready),         //     src20.ready
		.src20_valid         (cmd_xbar_demux_src20_valid),         //          .valid
		.src20_data          (cmd_xbar_demux_src20_data),          //          .data
		.src20_channel       (cmd_xbar_demux_src20_channel),       //          .channel
		.src20_startofpacket (cmd_xbar_demux_src20_startofpacket), //          .startofpacket
		.src20_endofpacket   (cmd_xbar_demux_src20_endofpacket),   //          .endofpacket
		.src21_ready         (cmd_xbar_demux_src21_ready),         //     src21.ready
		.src21_valid         (cmd_xbar_demux_src21_valid),         //          .valid
		.src21_data          (cmd_xbar_demux_src21_data),          //          .data
		.src21_channel       (cmd_xbar_demux_src21_channel),       //          .channel
		.src21_startofpacket (cmd_xbar_demux_src21_startofpacket), //          .startofpacket
		.src21_endofpacket   (cmd_xbar_demux_src21_endofpacket),   //          .endofpacket
		.src22_ready         (cmd_xbar_demux_src22_ready),         //     src22.ready
		.src22_valid         (cmd_xbar_demux_src22_valid),         //          .valid
		.src22_data          (cmd_xbar_demux_src22_data),          //          .data
		.src22_channel       (cmd_xbar_demux_src22_channel),       //          .channel
		.src22_startofpacket (cmd_xbar_demux_src22_startofpacket), //          .startofpacket
		.src22_endofpacket   (cmd_xbar_demux_src22_endofpacket),   //          .endofpacket
		.src23_ready         (cmd_xbar_demux_src23_ready),         //     src23.ready
		.src23_valid         (cmd_xbar_demux_src23_valid),         //          .valid
		.src23_data          (cmd_xbar_demux_src23_data),          //          .data
		.src23_channel       (cmd_xbar_demux_src23_channel),       //          .channel
		.src23_startofpacket (cmd_xbar_demux_src23_startofpacket), //          .startofpacket
		.src23_endofpacket   (cmd_xbar_demux_src23_endofpacket),   //          .endofpacket
		.src24_ready         (cmd_xbar_demux_src24_ready),         //     src24.ready
		.src24_valid         (cmd_xbar_demux_src24_valid),         //          .valid
		.src24_data          (cmd_xbar_demux_src24_data),          //          .data
		.src24_channel       (cmd_xbar_demux_src24_channel),       //          .channel
		.src24_startofpacket (cmd_xbar_demux_src24_startofpacket), //          .startofpacket
		.src24_endofpacket   (cmd_xbar_demux_src24_endofpacket)    //          .endofpacket
	);

	DE2_QSYS_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                (cpu_clk_for_sdram_clk),                 //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_001_src_ready),             //      sink.ready
		.sink_channel       (addr_router_001_src_channel),           //          .channel
		.sink_data          (addr_router_001_src_data),              //          .data
		.sink_startofpacket (addr_router_001_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_001_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_001_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	DE2_QSYS_cmd_xbar_demux_002 cmd_xbar_demux_002 (
		.clk                (clk_clk),                                //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),     // clk_reset.reset
		.sink_ready         (limiter_pipeline_source0_ready),         //      sink.ready
		.sink_channel       (limiter_pipeline_source0_channel),       //          .channel
		.sink_data          (limiter_pipeline_source0_data),          //          .data
		.sink_startofpacket (limiter_pipeline_source0_startofpacket), //          .startofpacket
		.sink_endofpacket   (limiter_pipeline_source0_endofpacket),   //          .endofpacket
		.sink_valid         (limiter_pipeline_source0_valid),         //          .valid
		.src0_ready         (cmd_xbar_demux_002_src0_ready),          //      src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),          //          .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),           //          .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),        //          .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket),    //          .endofpacket
		.src1_ready         (cmd_xbar_demux_002_src1_ready),          //      src1.ready
		.src1_valid         (cmd_xbar_demux_002_src1_valid),          //          .valid
		.src1_data          (cmd_xbar_demux_002_src1_data),           //          .data
		.src1_channel       (cmd_xbar_demux_002_src1_channel),        //          .channel
		.src1_startofpacket (cmd_xbar_demux_002_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_002_src1_endofpacket)     //          .endofpacket
	);

	DE2_QSYS_cmd_xbar_mux_006 cmd_xbar_mux_006 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_006_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_006_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_006_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_006_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_006_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_006_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src6_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src6_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src6_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src6_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src6_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src6_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	DE2_QSYS_cmd_xbar_mux_021 cmd_xbar_mux_021 (
		.clk                 (cpu_clk_for_sdram_clk),                 //       clk.clk
		.reset               (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_021_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_021_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_021_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_021_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_021_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_021_src_endofpacket),      //          .endofpacket
		.sink0_ready         (crosser_003_out_ready),                 //     sink0.ready
		.sink0_valid         (crosser_003_out_valid),                 //          .valid
		.sink0_channel       (crosser_003_out_channel),               //          .channel
		.sink0_data          (crosser_003_out_data),                  //          .data
		.sink0_startofpacket (crosser_003_out_startofpacket),         //          .startofpacket
		.sink0_endofpacket   (crosser_003_out_endofpacket),           //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (crosser_004_out_ready),                 //     sink2.ready
		.sink2_valid         (crosser_004_out_valid),                 //          .valid
		.sink2_channel       (crosser_004_out_channel),               //          .channel
		.sink2_data          (crosser_004_out_data),                  //          .data
		.sink2_startofpacket (crosser_004_out_startofpacket),         //          .startofpacket
		.sink2_endofpacket   (crosser_004_out_endofpacket)            //          .endofpacket
	);

	DE2_QSYS_cmd_xbar_demux_001 rsp_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket)    //          .endofpacket
	);

	DE2_QSYS_cmd_xbar_demux_001 rsp_xbar_demux_001 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	DE2_QSYS_cmd_xbar_demux_001 rsp_xbar_demux_002 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	DE2_QSYS_cmd_xbar_demux_001 rsp_xbar_demux_003 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	DE2_QSYS_cmd_xbar_demux_001 rsp_xbar_demux_004 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	DE2_QSYS_cmd_xbar_demux_001 rsp_xbar_demux_005 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	DE2_QSYS_cmd_xbar_demux_002 rsp_xbar_demux_006 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_006_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_006_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_006_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_006_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_006_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_006_src1_endofpacket)    //          .endofpacket
	);

	DE2_QSYS_cmd_xbar_demux_001 rsp_xbar_demux_007 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	DE2_QSYS_cmd_xbar_demux_001 rsp_xbar_demux_008 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	DE2_QSYS_cmd_xbar_demux_001 rsp_xbar_demux_009 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	DE2_QSYS_cmd_xbar_demux_001 rsp_xbar_demux_010 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	DE2_QSYS_cmd_xbar_demux_001 rsp_xbar_demux_011 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	DE2_QSYS_cmd_xbar_demux_001 rsp_xbar_demux_012 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	DE2_QSYS_cmd_xbar_demux_001 rsp_xbar_demux_013 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket)    //          .endofpacket
	);

	DE2_QSYS_cmd_xbar_demux_001 rsp_xbar_demux_014 (
		.clk                (clk_25_in_clk),                         //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_014_src_ready),               //      sink.ready
		.sink_channel       (id_router_014_src_channel),             //          .channel
		.sink_data          (id_router_014_src_data),                //          .data
		.sink_startofpacket (id_router_014_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_014_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_014_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket)    //          .endofpacket
	);

	DE2_QSYS_cmd_xbar_demux_001 rsp_xbar_demux_015 (
		.clk                (clk_40_in_clk),                         //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_015_src_ready),               //      sink.ready
		.sink_channel       (id_router_015_src_channel),             //          .channel
		.sink_data          (id_router_015_src_data),                //          .data
		.sink_startofpacket (id_router_015_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_015_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_015_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_015_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_015_src0_endofpacket)    //          .endofpacket
	);

	DE2_QSYS_cmd_xbar_demux_001 rsp_xbar_demux_016 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_016_src_ready),               //      sink.ready
		.sink_channel       (id_router_016_src_channel),             //          .channel
		.sink_data          (id_router_016_src_data),                //          .data
		.sink_startofpacket (id_router_016_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_016_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_016_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_016_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_016_src0_endofpacket)    //          .endofpacket
	);

	DE2_QSYS_cmd_xbar_demux_001 rsp_xbar_demux_017 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_017_src_ready),               //      sink.ready
		.sink_channel       (id_router_017_src_channel),             //          .channel
		.sink_data          (id_router_017_src_data),                //          .data
		.sink_startofpacket (id_router_017_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_017_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_017_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_017_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_017_src0_endofpacket)    //          .endofpacket
	);

	DE2_QSYS_cmd_xbar_demux_001 rsp_xbar_demux_018 (
		.clk                (cpu_clk_for_sdram_clk),                 //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_018_src_ready),               //      sink.ready
		.sink_channel       (id_router_018_src_channel),             //          .channel
		.sink_data          (id_router_018_src_data),                //          .data
		.sink_startofpacket (id_router_018_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_018_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_018_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_018_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_018_src0_endofpacket)    //          .endofpacket
	);

	DE2_QSYS_cmd_xbar_demux_001 rsp_xbar_demux_019 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_019_src_ready),               //      sink.ready
		.sink_channel       (id_router_019_src_channel),             //          .channel
		.sink_data          (id_router_019_src_data),                //          .data
		.sink_startofpacket (id_router_019_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_019_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_019_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_019_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_019_src0_endofpacket)    //          .endofpacket
	);

	DE2_QSYS_cmd_xbar_demux_001 rsp_xbar_demux_020 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_020_src_ready),               //      sink.ready
		.sink_channel       (id_router_020_src_channel),             //          .channel
		.sink_data          (id_router_020_src_data),                //          .data
		.sink_startofpacket (id_router_020_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_020_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_020_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_020_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_020_src0_endofpacket)    //          .endofpacket
	);

	DE2_QSYS_rsp_xbar_demux_021 rsp_xbar_demux_021 (
		.clk                (cpu_clk_for_sdram_clk),                 //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (width_adapter_001_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_001_src_channel),         //          .channel
		.sink_data          (width_adapter_001_src_data),            //          .data
		.sink_startofpacket (width_adapter_001_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_001_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_001_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_021_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_021_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_021_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_021_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_021_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_021_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_021_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_021_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_021_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_021_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_021_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_021_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_021_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_021_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_021_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_021_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_021_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_021_src2_endofpacket)    //          .endofpacket
	);

	DE2_QSYS_cmd_xbar_demux_001 rsp_xbar_demux_022 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_022_src_ready),               //      sink.ready
		.sink_channel       (id_router_022_src_channel),             //          .channel
		.sink_data          (id_router_022_src_data),                //          .data
		.sink_startofpacket (id_router_022_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_022_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_022_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_022_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_022_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_022_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_022_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_022_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_022_src0_endofpacket)    //          .endofpacket
	);

	DE2_QSYS_cmd_xbar_demux_001 rsp_xbar_demux_023 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_023_src_ready),               //      sink.ready
		.sink_channel       (id_router_023_src_channel),             //          .channel
		.sink_data          (id_router_023_src_data),                //          .data
		.sink_startofpacket (id_router_023_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_023_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_023_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_023_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_023_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_023_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_023_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_023_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_023_src0_endofpacket)    //          .endofpacket
	);

	DE2_QSYS_cmd_xbar_demux_001 rsp_xbar_demux_024 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_024_src_ready),               //      sink.ready
		.sink_channel       (id_router_024_src_channel),             //          .channel
		.sink_data          (id_router_024_src_data),                //          .data
		.sink_startofpacket (id_router_024_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_024_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_024_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_024_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_024_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_024_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_024_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_024_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_024_src0_endofpacket)    //          .endofpacket
	);

	DE2_QSYS_rsp_xbar_mux rsp_xbar_mux (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready            (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid            (rsp_xbar_mux_src_valid),                //          .valid
		.src_data             (rsp_xbar_mux_src_data),                 //          .data
		.src_channel          (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket    (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_010_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_011_src0_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_012_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_013_src0_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.sink14_ready         (crosser_005_out_ready),                 //    sink14.ready
		.sink14_valid         (crosser_005_out_valid),                 //          .valid
		.sink14_channel       (crosser_005_out_channel),               //          .channel
		.sink14_data          (crosser_005_out_data),                  //          .data
		.sink14_startofpacket (crosser_005_out_startofpacket),         //          .startofpacket
		.sink14_endofpacket   (crosser_005_out_endofpacket),           //          .endofpacket
		.sink15_ready         (crosser_006_out_ready),                 //    sink15.ready
		.sink15_valid         (crosser_006_out_valid),                 //          .valid
		.sink15_channel       (crosser_006_out_channel),               //          .channel
		.sink15_data          (crosser_006_out_data),                  //          .data
		.sink15_startofpacket (crosser_006_out_startofpacket),         //          .startofpacket
		.sink15_endofpacket   (crosser_006_out_endofpacket),           //          .endofpacket
		.sink16_ready         (rsp_xbar_demux_016_src0_ready),         //    sink16.ready
		.sink16_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.sink16_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.sink16_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.sink16_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.sink16_endofpacket   (rsp_xbar_demux_016_src0_endofpacket),   //          .endofpacket
		.sink17_ready         (rsp_xbar_demux_017_src0_ready),         //    sink17.ready
		.sink17_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.sink17_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.sink17_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.sink17_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.sink17_endofpacket   (rsp_xbar_demux_017_src0_endofpacket),   //          .endofpacket
		.sink18_ready         (crosser_007_out_ready),                 //    sink18.ready
		.sink18_valid         (crosser_007_out_valid),                 //          .valid
		.sink18_channel       (crosser_007_out_channel),               //          .channel
		.sink18_data          (crosser_007_out_data),                  //          .data
		.sink18_startofpacket (crosser_007_out_startofpacket),         //          .startofpacket
		.sink18_endofpacket   (crosser_007_out_endofpacket),           //          .endofpacket
		.sink19_ready         (rsp_xbar_demux_019_src0_ready),         //    sink19.ready
		.sink19_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.sink19_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.sink19_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.sink19_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.sink19_endofpacket   (rsp_xbar_demux_019_src0_endofpacket),   //          .endofpacket
		.sink20_ready         (rsp_xbar_demux_020_src0_ready),         //    sink20.ready
		.sink20_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.sink20_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.sink20_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.sink20_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.sink20_endofpacket   (rsp_xbar_demux_020_src0_endofpacket),   //          .endofpacket
		.sink21_ready         (crosser_008_out_ready),                 //    sink21.ready
		.sink21_valid         (crosser_008_out_valid),                 //          .valid
		.sink21_channel       (crosser_008_out_channel),               //          .channel
		.sink21_data          (crosser_008_out_data),                  //          .data
		.sink21_startofpacket (crosser_008_out_startofpacket),         //          .startofpacket
		.sink21_endofpacket   (crosser_008_out_endofpacket),           //          .endofpacket
		.sink22_ready         (rsp_xbar_demux_022_src0_ready),         //    sink22.ready
		.sink22_valid         (rsp_xbar_demux_022_src0_valid),         //          .valid
		.sink22_channel       (rsp_xbar_demux_022_src0_channel),       //          .channel
		.sink22_data          (rsp_xbar_demux_022_src0_data),          //          .data
		.sink22_startofpacket (rsp_xbar_demux_022_src0_startofpacket), //          .startofpacket
		.sink22_endofpacket   (rsp_xbar_demux_022_src0_endofpacket),   //          .endofpacket
		.sink23_ready         (rsp_xbar_demux_023_src0_ready),         //    sink23.ready
		.sink23_valid         (rsp_xbar_demux_023_src0_valid),         //          .valid
		.sink23_channel       (rsp_xbar_demux_023_src0_channel),       //          .channel
		.sink23_data          (rsp_xbar_demux_023_src0_data),          //          .data
		.sink23_startofpacket (rsp_xbar_demux_023_src0_startofpacket), //          .startofpacket
		.sink23_endofpacket   (rsp_xbar_demux_023_src0_endofpacket),   //          .endofpacket
		.sink24_ready         (rsp_xbar_demux_024_src0_ready),         //    sink24.ready
		.sink24_valid         (rsp_xbar_demux_024_src0_valid),         //          .valid
		.sink24_channel       (rsp_xbar_demux_024_src0_channel),       //          .channel
		.sink24_data          (rsp_xbar_demux_024_src0_data),          //          .data
		.sink24_startofpacket (rsp_xbar_demux_024_src0_startofpacket), //          .startofpacket
		.sink24_endofpacket   (rsp_xbar_demux_024_src0_endofpacket)    //          .endofpacket
	);

	DE2_QSYS_rsp_xbar_mux_002 rsp_xbar_mux_002 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_002_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_002_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_006_src1_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_006_src1_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_006_src1_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_006_src1_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_006_src1_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_006_src1_endofpacket),   //          .endofpacket
		.sink1_ready         (crosser_009_out_ready),                 //     sink1.ready
		.sink1_valid         (crosser_009_out_valid),                 //          .valid
		.sink1_channel       (crosser_009_out_channel),               //          .channel
		.sink1_data          (crosser_009_out_data),                  //          .data
		.sink1_startofpacket (crosser_009_out_startofpacket),         //          .startofpacket
		.sink1_endofpacket   (crosser_009_out_endofpacket)            //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (81),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (84),
		.IN_PKT_BURSTWRAP_L            (82),
		.IN_PKT_BURST_SIZE_H           (87),
		.IN_PKT_BURST_SIZE_L           (85),
		.IN_PKT_RESPONSE_STATUS_H      (113),
		.IN_PKT_RESPONSE_STATUS_L      (112),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (89),
		.IN_PKT_BURST_TYPE_L           (88),
		.IN_ST_DATA_W                  (114),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (63),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (69),
		.OUT_PKT_BURST_SIZE_L          (67),
		.OUT_PKT_RESPONSE_STATUS_H     (95),
		.OUT_PKT_RESPONSE_STATUS_L     (94),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (71),
		.OUT_PKT_BURST_TYPE_L          (70),
		.OUT_ST_DATA_W                 (96),
		.ST_CHANNEL_W                  (25),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter (
		.clk                  (cpu_clk_for_sdram_clk),              //       clk.clk
		.reset                (rst_controller_004_reset_out_reset), // clk_reset.reset
		.in_valid             (cmd_xbar_mux_021_src_valid),         //      sink.valid
		.in_channel           (cmd_xbar_mux_021_src_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_mux_021_src_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_mux_021_src_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_mux_021_src_ready),         //          .ready
		.in_data              (cmd_xbar_mux_021_src_data),          //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_src_data),             //          .data
		.out_channel          (width_adapter_src_channel),          //          .channel
		.out_valid            (width_adapter_src_valid),            //          .valid
		.out_ready            (width_adapter_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                              // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (63),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (66),
		.IN_PKT_BURSTWRAP_L            (64),
		.IN_PKT_BURST_SIZE_H           (69),
		.IN_PKT_BURST_SIZE_L           (67),
		.IN_PKT_RESPONSE_STATUS_H      (95),
		.IN_PKT_RESPONSE_STATUS_L      (94),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (71),
		.IN_PKT_BURST_TYPE_L           (70),
		.IN_ST_DATA_W                  (96),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (81),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (87),
		.OUT_PKT_BURST_SIZE_L          (85),
		.OUT_PKT_RESPONSE_STATUS_H     (113),
		.OUT_PKT_RESPONSE_STATUS_L     (112),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (89),
		.OUT_PKT_BURST_TYPE_L          (88),
		.OUT_ST_DATA_W                 (114),
		.ST_CHANNEL_W                  (25),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (1)
	) width_adapter_001 (
		.clk                  (cpu_clk_for_sdram_clk),               //       clk.clk
		.reset                (rst_controller_004_reset_out_reset),  // clk_reset.reset
		.in_valid             (id_router_021_src_valid),             //      sink.valid
		.in_channel           (id_router_021_src_channel),           //          .channel
		.in_startofpacket     (id_router_021_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_021_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_021_src_ready),             //          .ready
		.in_data              (id_router_021_src_data),              //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_001_src_data),          //          .data
		.out_channel          (width_adapter_001_src_channel),       //          .channel
		.out_valid            (width_adapter_001_src_valid),         //          .valid
		.out_ready            (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (114),
		.BITS_PER_SYMBOL     (114),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (25),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser (
		.in_clk            (clk_clk),                            //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset), //  in_clk_reset.reset
		.out_clk           (clk_25_in_clk),                      //       out_clk.clk
		.out_reset         (rst_controller_002_reset_out_reset), // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_src14_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_src14_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_src14_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src14_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_src14_channel),       //              .channel
		.in_data           (cmd_xbar_demux_src14_data),          //              .data
		.out_ready         (crosser_out_ready),                  //           out.ready
		.out_valid         (crosser_out_valid),                  //              .valid
		.out_startofpacket (crosser_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_out_channel),                //              .channel
		.out_data          (crosser_out_data),                   //              .data
		.in_empty          (1'b0),                               //   (terminated)
		.in_error          (1'b0),                               //   (terminated)
		.out_empty         (),                                   //   (terminated)
		.out_error         ()                                    //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (114),
		.BITS_PER_SYMBOL     (114),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (25),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_001 (
		.in_clk            (clk_clk),                            //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset), //  in_clk_reset.reset
		.out_clk           (clk_40_in_clk),                      //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset), // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_src15_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_src15_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_src15_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src15_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_src15_channel),       //              .channel
		.in_data           (cmd_xbar_demux_src15_data),          //              .data
		.out_ready         (crosser_001_out_ready),              //           out.ready
		.out_valid         (crosser_001_out_valid),              //              .valid
		.out_startofpacket (crosser_001_out_startofpacket),      //              .startofpacket
		.out_endofpacket   (crosser_001_out_endofpacket),        //              .endofpacket
		.out_channel       (crosser_001_out_channel),            //              .channel
		.out_data          (crosser_001_out_data),               //              .data
		.in_empty          (1'b0),                               //   (terminated)
		.in_error          (1'b0),                               //   (terminated)
		.out_empty         (),                                   //   (terminated)
		.out_error         ()                                    //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (114),
		.BITS_PER_SYMBOL     (114),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (25),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_002 (
		.in_clk            (clk_clk),                            //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset), //  in_clk_reset.reset
		.out_clk           (cpu_clk_for_sdram_clk),              //       out_clk.clk
		.out_reset         (rst_controller_004_reset_out_reset), // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_src18_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_src18_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_src18_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src18_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_src18_channel),       //              .channel
		.in_data           (cmd_xbar_demux_src18_data),          //              .data
		.out_ready         (crosser_002_out_ready),              //           out.ready
		.out_valid         (crosser_002_out_valid),              //              .valid
		.out_startofpacket (crosser_002_out_startofpacket),      //              .startofpacket
		.out_endofpacket   (crosser_002_out_endofpacket),        //              .endofpacket
		.out_channel       (crosser_002_out_channel),            //              .channel
		.out_data          (crosser_002_out_data),               //              .data
		.in_empty          (1'b0),                               //   (terminated)
		.in_error          (1'b0),                               //   (terminated)
		.out_empty         (),                                   //   (terminated)
		.out_error         ()                                    //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (114),
		.BITS_PER_SYMBOL     (114),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (25),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_003 (
		.in_clk            (clk_clk),                            //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset), //  in_clk_reset.reset
		.out_clk           (cpu_clk_for_sdram_clk),              //       out_clk.clk
		.out_reset         (rst_controller_004_reset_out_reset), // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_src21_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_src21_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_src21_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src21_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_src21_channel),       //              .channel
		.in_data           (cmd_xbar_demux_src21_data),          //              .data
		.out_ready         (crosser_003_out_ready),              //           out.ready
		.out_valid         (crosser_003_out_valid),              //              .valid
		.out_startofpacket (crosser_003_out_startofpacket),      //              .startofpacket
		.out_endofpacket   (crosser_003_out_endofpacket),        //              .endofpacket
		.out_channel       (crosser_003_out_channel),            //              .channel
		.out_data          (crosser_003_out_data),               //              .data
		.in_empty          (1'b0),                               //   (terminated)
		.in_error          (1'b0),                               //   (terminated)
		.out_empty         (),                                   //   (terminated)
		.out_error         ()                                    //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (114),
		.BITS_PER_SYMBOL     (114),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (25),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_004 (
		.in_clk            (clk_clk),                               //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (cpu_clk_for_sdram_clk),                 //       out_clk.clk
		.out_reset         (rst_controller_004_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_002_src1_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_002_src1_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_002_src1_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_002_src1_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_002_src1_channel),       //              .channel
		.in_data           (cmd_xbar_demux_002_src1_data),          //              .data
		.out_ready         (crosser_004_out_ready),                 //           out.ready
		.out_valid         (crosser_004_out_valid),                 //              .valid
		.out_startofpacket (crosser_004_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_004_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_004_out_channel),               //              .channel
		.out_data          (crosser_004_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (114),
		.BITS_PER_SYMBOL     (114),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (25),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_005 (
		.in_clk            (clk_25_in_clk),                         //        in_clk.clk
		.in_reset          (rst_controller_002_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (clk_clk),                               //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_014_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_014_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_014_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_014_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_014_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_014_src0_data),          //              .data
		.out_ready         (crosser_005_out_ready),                 //           out.ready
		.out_valid         (crosser_005_out_valid),                 //              .valid
		.out_startofpacket (crosser_005_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_005_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_005_out_channel),               //              .channel
		.out_data          (crosser_005_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (114),
		.BITS_PER_SYMBOL     (114),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (25),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_006 (
		.in_clk            (clk_40_in_clk),                         //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (clk_clk),                               //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_015_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_015_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_015_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_015_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_015_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_015_src0_data),          //              .data
		.out_ready         (crosser_006_out_ready),                 //           out.ready
		.out_valid         (crosser_006_out_valid),                 //              .valid
		.out_startofpacket (crosser_006_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_006_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_006_out_channel),               //              .channel
		.out_data          (crosser_006_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (114),
		.BITS_PER_SYMBOL     (114),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (25),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_007 (
		.in_clk            (cpu_clk_for_sdram_clk),                 //        in_clk.clk
		.in_reset          (rst_controller_004_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (clk_clk),                               //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_018_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_018_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_018_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_018_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_018_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_018_src0_data),          //              .data
		.out_ready         (crosser_007_out_ready),                 //           out.ready
		.out_valid         (crosser_007_out_valid),                 //              .valid
		.out_startofpacket (crosser_007_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_007_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_007_out_channel),               //              .channel
		.out_data          (crosser_007_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (114),
		.BITS_PER_SYMBOL     (114),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (25),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_008 (
		.in_clk            (cpu_clk_for_sdram_clk),                 //        in_clk.clk
		.in_reset          (rst_controller_004_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (clk_clk),                               //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_021_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_021_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_021_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_021_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_021_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_021_src0_data),          //              .data
		.out_ready         (crosser_008_out_ready),                 //           out.ready
		.out_valid         (crosser_008_out_valid),                 //              .valid
		.out_startofpacket (crosser_008_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_008_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_008_out_channel),               //              .channel
		.out_data          (crosser_008_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (114),
		.BITS_PER_SYMBOL     (114),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (25),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_009 (
		.in_clk            (cpu_clk_for_sdram_clk),                 //        in_clk.clk
		.in_reset          (rst_controller_004_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (clk_clk),                               //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_021_src2_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_021_src2_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_021_src2_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_021_src2_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_021_src2_channel),       //              .channel
		.in_data           (rsp_xbar_demux_021_src2_data),          //              .data
		.out_ready         (crosser_009_out_ready),                 //           out.ready
		.out_valid         (crosser_009_out_valid),                 //              .valid
		.out_startofpacket (crosser_009_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_009_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_009_out_channel),               //              .channel
		.out_data          (crosser_009_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (25),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) limiter_pipeline (
		.clk               (clk_clk),                                //       cr0.clk
		.reset             (rst_controller_001_reset_out_reset),     // cr0_reset.reset
		.in_ready          (limiter_cmd_src_ready),                  //     sink0.ready
		.in_valid          (limiter_cmd_src_valid),                  //          .valid
		.in_startofpacket  (limiter_cmd_src_startofpacket),          //          .startofpacket
		.in_endofpacket    (limiter_cmd_src_endofpacket),            //          .endofpacket
		.in_data           (limiter_cmd_src_data),                   //          .data
		.in_channel        (limiter_cmd_src_channel),                //          .channel
		.out_ready         (limiter_pipeline_source0_ready),         //   source0.ready
		.out_valid         (limiter_pipeline_source0_valid),         //          .valid
		.out_startofpacket (limiter_pipeline_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (limiter_pipeline_source0_endofpacket),   //          .endofpacket
		.out_data          (limiter_pipeline_source0_data),          //          .data
		.out_channel       (limiter_pipeline_source0_channel),       //          .channel
		.in_empty          (1'b0),                                   // (terminated)
		.out_empty         (),                                       // (terminated)
		.out_error         (),                                       // (terminated)
		.in_error          (1'b0)                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (25),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) limiter_pipeline_001 (
		.clk               (clk_clk),                                    //       cr0.clk
		.reset             (rst_controller_001_reset_out_reset),         // cr0_reset.reset
		.in_ready          (rsp_xbar_mux_002_src_ready),                 //     sink0.ready
		.in_valid          (rsp_xbar_mux_002_src_valid),                 //          .valid
		.in_startofpacket  (rsp_xbar_mux_002_src_startofpacket),         //          .startofpacket
		.in_endofpacket    (rsp_xbar_mux_002_src_endofpacket),           //          .endofpacket
		.in_data           (rsp_xbar_mux_002_src_data),                  //          .data
		.in_channel        (rsp_xbar_mux_002_src_channel),               //          .channel
		.out_ready         (limiter_pipeline_001_source0_ready),         //   source0.ready
		.out_valid         (limiter_pipeline_001_source0_valid),         //          .valid
		.out_startofpacket (limiter_pipeline_001_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (limiter_pipeline_001_source0_endofpacket),   //          .endofpacket
		.out_data          (limiter_pipeline_001_source0_data),          //          .data
		.out_channel       (limiter_pipeline_001_source0_channel),       //          .channel
		.in_empty          (1'b0),                                       // (terminated)
		.out_empty         (),                                           // (terminated)
		.out_error         (),                                           // (terminated)
		.in_error          (1'b0)                                        // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (25),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline (
		.clk               (clk_clk),                              //       cr0.clk
		.reset             (rst_controller_reset_out_reset),       // cr0_reset.reset
		.in_ready          (cmd_xbar_demux_src0_ready),            //     sink0.ready
		.in_valid          (cmd_xbar_demux_src0_valid),            //          .valid
		.in_startofpacket  (cmd_xbar_demux_src0_startofpacket),    //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src0_endofpacket),      //          .endofpacket
		.in_data           (cmd_xbar_demux_src0_data),             //          .data
		.in_channel        (cmd_xbar_demux_src0_channel),          //          .channel
		.out_ready         (agent_pipeline_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_source0_data),          //          .data
		.out_channel       (agent_pipeline_source0_channel),       //          .channel
		.in_empty          (1'b0),                                 // (terminated)
		.out_empty         (),                                     // (terminated)
		.out_error         (),                                     // (terminated)
		.in_error          (1'b0)                                  // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_001 (
		.clk               (clk_clk),                                                                                //       cr0.clk
		.reset             (rst_controller_reset_out_reset),                                                         // cr0_reset.reset
		.in_ready          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_001_source0_ready),                                                       //   source0.ready
		.out_valid         (agent_pipeline_001_source0_valid),                                                       //          .valid
		.out_startofpacket (agent_pipeline_001_source0_startofpacket),                                               //          .startofpacket
		.out_endofpacket   (agent_pipeline_001_source0_endofpacket),                                                 //          .endofpacket
		.out_data          (agent_pipeline_001_source0_data),                                                        //          .data
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_channel       (),                                                                                       // (terminated)
		.in_channel        (1'b0)                                                                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (25),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_002 (
		.clk               (clk_clk),                                  //       cr0.clk
		.reset             (rst_controller_reset_out_reset),           // cr0_reset.reset
		.in_ready          (cmd_xbar_demux_src1_ready),                //     sink0.ready
		.in_valid          (cmd_xbar_demux_src1_valid),                //          .valid
		.in_startofpacket  (cmd_xbar_demux_src1_startofpacket),        //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src1_endofpacket),          //          .endofpacket
		.in_data           (cmd_xbar_demux_src1_data),                 //          .data
		.in_channel        (cmd_xbar_demux_src1_channel),              //          .channel
		.out_ready         (agent_pipeline_002_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_002_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_002_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_002_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_002_source0_data),          //          .data
		.out_channel       (agent_pipeline_002_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_003 (
		.clk               (clk_clk),                                                                             //       cr0.clk
		.reset             (rst_controller_reset_out_reset),                                                      // cr0_reset.reset
		.in_ready          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_003_source0_ready),                                                    //   source0.ready
		.out_valid         (agent_pipeline_003_source0_valid),                                                    //          .valid
		.out_startofpacket (agent_pipeline_003_source0_startofpacket),                                            //          .startofpacket
		.out_endofpacket   (agent_pipeline_003_source0_endofpacket),                                              //          .endofpacket
		.out_data          (agent_pipeline_003_source0_data),                                                     //          .data
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_channel       (),                                                                                    // (terminated)
		.in_channel        (1'b0)                                                                                 // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (25),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_004 (
		.clk               (clk_clk),                                  //       cr0.clk
		.reset             (rst_controller_reset_out_reset),           // cr0_reset.reset
		.in_ready          (cmd_xbar_demux_src2_ready),                //     sink0.ready
		.in_valid          (cmd_xbar_demux_src2_valid),                //          .valid
		.in_startofpacket  (cmd_xbar_demux_src2_startofpacket),        //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src2_endofpacket),          //          .endofpacket
		.in_data           (cmd_xbar_demux_src2_data),                 //          .data
		.in_channel        (cmd_xbar_demux_src2_channel),              //          .channel
		.out_ready         (agent_pipeline_004_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_004_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_004_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_004_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_004_source0_data),          //          .data
		.out_channel       (agent_pipeline_004_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_005 (
		.clk               (clk_clk),                                                                         //       cr0.clk
		.reset             (rst_controller_reset_out_reset),                                                  // cr0_reset.reset
		.in_ready          (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (audio_data_fregen_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_005_source0_ready),                                                //   source0.ready
		.out_valid         (agent_pipeline_005_source0_valid),                                                //          .valid
		.out_startofpacket (agent_pipeline_005_source0_startofpacket),                                        //          .startofpacket
		.out_endofpacket   (agent_pipeline_005_source0_endofpacket),                                          //          .endofpacket
		.out_data          (agent_pipeline_005_source0_data),                                                 //          .data
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_channel       (),                                                                                // (terminated)
		.in_channel        (1'b0)                                                                             // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (25),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_006 (
		.clk               (clk_clk),                                  //       cr0.clk
		.reset             (rst_controller_reset_out_reset),           // cr0_reset.reset
		.in_ready          (cmd_xbar_demux_src3_ready),                //     sink0.ready
		.in_valid          (cmd_xbar_demux_src3_valid),                //          .valid
		.in_startofpacket  (cmd_xbar_demux_src3_startofpacket),        //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src3_endofpacket),          //          .endofpacket
		.in_data           (cmd_xbar_demux_src3_data),                 //          .data
		.in_channel        (cmd_xbar_demux_src3_channel),              //          .channel
		.out_ready         (agent_pipeline_006_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_006_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_006_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_006_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_006_source0_data),          //          .data
		.out_channel       (agent_pipeline_006_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_007 (
		.clk               (clk_clk),                                                                   //       cr0.clk
		.reset             (rst_controller_reset_out_reset),                                            // cr0_reset.reset
		.in_ready          (audio_empty_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (audio_empty_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (audio_empty_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (audio_empty_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (audio_empty_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_007_source0_ready),                                          //   source0.ready
		.out_valid         (agent_pipeline_007_source0_valid),                                          //          .valid
		.out_startofpacket (agent_pipeline_007_source0_startofpacket),                                  //          .startofpacket
		.out_endofpacket   (agent_pipeline_007_source0_endofpacket),                                    //          .endofpacket
		.out_data          (agent_pipeline_007_source0_data),                                           //          .data
		.in_empty          (1'b0),                                                                      // (terminated)
		.out_empty         (),                                                                          // (terminated)
		.out_error         (),                                                                          // (terminated)
		.in_error          (1'b0),                                                                      // (terminated)
		.out_channel       (),                                                                          // (terminated)
		.in_channel        (1'b0)                                                                       // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (25),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_008 (
		.clk               (clk_clk),                                  //       cr0.clk
		.reset             (rst_controller_reset_out_reset),           // cr0_reset.reset
		.in_ready          (cmd_xbar_demux_src4_ready),                //     sink0.ready
		.in_valid          (cmd_xbar_demux_src4_valid),                //          .valid
		.in_startofpacket  (cmd_xbar_demux_src4_startofpacket),        //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src4_endofpacket),          //          .endofpacket
		.in_data           (cmd_xbar_demux_src4_data),                 //          .data
		.in_channel        (cmd_xbar_demux_src4_channel),              //          .channel
		.out_ready         (agent_pipeline_008_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_008_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_008_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_008_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_008_source0_data),          //          .data
		.out_channel       (agent_pipeline_008_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_009 (
		.clk               (clk_clk),                                                                       //       cr0.clk
		.reset             (rst_controller_reset_out_reset),                                                // cr0_reset.reset
		.in_ready          (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (audio_fifo_full_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_009_source0_ready),                                              //   source0.ready
		.out_valid         (agent_pipeline_009_source0_valid),                                              //          .valid
		.out_startofpacket (agent_pipeline_009_source0_startofpacket),                                      //          .startofpacket
		.out_endofpacket   (agent_pipeline_009_source0_endofpacket),                                        //          .endofpacket
		.out_data          (agent_pipeline_009_source0_data),                                               //          .data
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_channel       (),                                                                              // (terminated)
		.in_channel        (1'b0)                                                                           // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (25),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_010 (
		.clk               (clk_clk),                                  //       cr0.clk
		.reset             (rst_controller_reset_out_reset),           // cr0_reset.reset
		.in_ready          (cmd_xbar_demux_src5_ready),                //     sink0.ready
		.in_valid          (cmd_xbar_demux_src5_valid),                //          .valid
		.in_startofpacket  (cmd_xbar_demux_src5_startofpacket),        //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src5_endofpacket),          //          .endofpacket
		.in_data           (cmd_xbar_demux_src5_data),                 //          .data
		.in_channel        (cmd_xbar_demux_src5_channel),              //          .channel
		.out_ready         (agent_pipeline_010_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_010_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_010_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_010_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_010_source0_data),          //          .data
		.out_channel       (agent_pipeline_010_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_011 (
		.clk               (clk_clk),                                                                       //       cr0.clk
		.reset             (rst_controller_reset_out_reset),                                                // cr0_reset.reset
		.in_ready          (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (audio_fifo_used_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_011_source0_ready),                                              //   source0.ready
		.out_valid         (agent_pipeline_011_source0_valid),                                              //          .valid
		.out_startofpacket (agent_pipeline_011_source0_startofpacket),                                      //          .startofpacket
		.out_endofpacket   (agent_pipeline_011_source0_endofpacket),                                        //          .endofpacket
		.out_data          (agent_pipeline_011_source0_data),                                               //          .data
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_channel       (),                                                                              // (terminated)
		.in_channel        (1'b0)                                                                           // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (25),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_012 (
		.clk               (clk_clk),                                  //       cr0.clk
		.reset             (rst_controller_001_reset_out_reset),       // cr0_reset.reset
		.in_ready          (cmd_xbar_mux_006_src_ready),               //     sink0.ready
		.in_valid          (cmd_xbar_mux_006_src_valid),               //          .valid
		.in_startofpacket  (cmd_xbar_mux_006_src_startofpacket),       //          .startofpacket
		.in_endofpacket    (cmd_xbar_mux_006_src_endofpacket),         //          .endofpacket
		.in_data           (cmd_xbar_mux_006_src_data),                //          .data
		.in_channel        (cmd_xbar_mux_006_src_channel),             //          .channel
		.out_ready         (agent_pipeline_012_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_012_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_012_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_012_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_012_source0_data),          //          .data
		.out_channel       (agent_pipeline_012_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_013 (
		.clk               (clk_clk),                                                                          //       cr0.clk
		.reset             (rst_controller_001_reset_out_reset),                                               // cr0_reset.reset
		.in_ready          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_013_source0_ready),                                                 //   source0.ready
		.out_valid         (agent_pipeline_013_source0_valid),                                                 //          .valid
		.out_startofpacket (agent_pipeline_013_source0_startofpacket),                                         //          .startofpacket
		.out_endofpacket   (agent_pipeline_013_source0_endofpacket),                                           //          .endofpacket
		.out_data          (agent_pipeline_013_source0_data),                                                  //          .data
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_channel       (),                                                                                 // (terminated)
		.in_channel        (1'b0)                                                                              // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (25),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_014 (
		.clk               (clk_clk),                                  //       cr0.clk
		.reset             (rst_controller_reset_out_reset),           // cr0_reset.reset
		.in_ready          (cmd_xbar_demux_src7_ready),                //     sink0.ready
		.in_valid          (cmd_xbar_demux_src7_valid),                //          .valid
		.in_startofpacket  (cmd_xbar_demux_src7_startofpacket),        //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src7_endofpacket),          //          .endofpacket
		.in_data           (cmd_xbar_demux_src7_data),                 //          .data
		.in_channel        (cmd_xbar_demux_src7_channel),              //          .channel
		.out_ready         (agent_pipeline_014_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_014_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_014_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_014_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_014_source0_data),          //          .data
		.out_channel       (agent_pipeline_014_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_015 (
		.clk               (clk_clk),                                                                            //       cr0.clk
		.reset             (rst_controller_reset_out_reset),                                                     // cr0_reset.reset
		.in_ready          (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (audio_out_data_audio_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_015_source0_ready),                                                   //   source0.ready
		.out_valid         (agent_pipeline_015_source0_valid),                                                   //          .valid
		.out_startofpacket (agent_pipeline_015_source0_startofpacket),                                           //          .startofpacket
		.out_endofpacket   (agent_pipeline_015_source0_endofpacket),                                             //          .endofpacket
		.out_data          (agent_pipeline_015_source0_data),                                                    //          .data
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_channel       (),                                                                                   // (terminated)
		.in_channel        (1'b0)                                                                                // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (25),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_016 (
		.clk               (clk_clk),                                  //       cr0.clk
		.reset             (rst_controller_reset_out_reset),           // cr0_reset.reset
		.in_ready          (cmd_xbar_demux_src8_ready),                //     sink0.ready
		.in_valid          (cmd_xbar_demux_src8_valid),                //          .valid
		.in_startofpacket  (cmd_xbar_demux_src8_startofpacket),        //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src8_endofpacket),          //          .endofpacket
		.in_data           (cmd_xbar_demux_src8_data),                 //          .data
		.in_channel        (cmd_xbar_demux_src8_channel),              //          .channel
		.out_ready         (agent_pipeline_016_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_016_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_016_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_016_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_016_source0_data),          //          .data
		.out_channel       (agent_pipeline_016_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_017 (
		.clk               (clk_clk),                                                                       //       cr0.clk
		.reset             (rst_controller_reset_out_reset),                                                // cr0_reset.reset
		.in_ready          (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (audio_out_pause_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_017_source0_ready),                                              //   source0.ready
		.out_valid         (agent_pipeline_017_source0_valid),                                              //          .valid
		.out_startofpacket (agent_pipeline_017_source0_startofpacket),                                      //          .startofpacket
		.out_endofpacket   (agent_pipeline_017_source0_endofpacket),                                        //          .endofpacket
		.out_data          (agent_pipeline_017_source0_data),                                               //          .data
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_channel       (),                                                                              // (terminated)
		.in_channel        (1'b0)                                                                           // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (25),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_018 (
		.clk               (clk_clk),                                  //       cr0.clk
		.reset             (rst_controller_reset_out_reset),           // cr0_reset.reset
		.in_ready          (cmd_xbar_demux_src9_ready),                //     sink0.ready
		.in_valid          (cmd_xbar_demux_src9_valid),                //          .valid
		.in_startofpacket  (cmd_xbar_demux_src9_startofpacket),        //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src9_endofpacket),          //          .endofpacket
		.in_data           (cmd_xbar_demux_src9_data),                 //          .data
		.in_channel        (cmd_xbar_demux_src9_channel),              //          .channel
		.out_ready         (agent_pipeline_018_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_018_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_018_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_018_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_018_source0_data),          //          .data
		.out_channel       (agent_pipeline_018_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_019 (
		.clk               (clk_clk),                                                                      //       cr0.clk
		.reset             (rst_controller_reset_out_reset),                                               // cr0_reset.reset
		.in_ready          (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (audio_out_stop_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_019_source0_ready),                                             //   source0.ready
		.out_valid         (agent_pipeline_019_source0_valid),                                             //          .valid
		.out_startofpacket (agent_pipeline_019_source0_startofpacket),                                     //          .startofpacket
		.out_endofpacket   (agent_pipeline_019_source0_endofpacket),                                       //          .endofpacket
		.out_data          (agent_pipeline_019_source0_data),                                              //          .data
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_channel       (),                                                                             // (terminated)
		.in_channel        (1'b0)                                                                          // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (25),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_020 (
		.clk               (clk_clk),                                  //       cr0.clk
		.reset             (rst_controller_reset_out_reset),           // cr0_reset.reset
		.in_ready          (cmd_xbar_demux_src10_ready),               //     sink0.ready
		.in_valid          (cmd_xbar_demux_src10_valid),               //          .valid
		.in_startofpacket  (cmd_xbar_demux_src10_startofpacket),       //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src10_endofpacket),         //          .endofpacket
		.in_data           (cmd_xbar_demux_src10_data),                //          .data
		.in_channel        (cmd_xbar_demux_src10_channel),             //          .channel
		.out_ready         (agent_pipeline_020_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_020_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_020_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_020_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_020_source0_data),          //          .data
		.out_channel       (agent_pipeline_020_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_021 (
		.clk               (clk_clk),                                                             //       cr0.clk
		.reset             (rst_controller_reset_out_reset),                                      // cr0_reset.reset
		.in_ready          (timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (timer_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_021_source0_ready),                                    //   source0.ready
		.out_valid         (agent_pipeline_021_source0_valid),                                    //          .valid
		.out_startofpacket (agent_pipeline_021_source0_startofpacket),                            //          .startofpacket
		.out_endofpacket   (agent_pipeline_021_source0_endofpacket),                              //          .endofpacket
		.out_data          (agent_pipeline_021_source0_data),                                     //          .data
		.in_empty          (1'b0),                                                                // (terminated)
		.out_empty         (),                                                                    // (terminated)
		.out_error         (),                                                                    // (terminated)
		.in_error          (1'b0),                                                                // (terminated)
		.out_channel       (),                                                                    // (terminated)
		.in_channel        (1'b0)                                                                 // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (25),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_022 (
		.clk               (clk_clk),                                  //       cr0.clk
		.reset             (rst_controller_reset_out_reset),           // cr0_reset.reset
		.in_ready          (cmd_xbar_demux_src11_ready),               //     sink0.ready
		.in_valid          (cmd_xbar_demux_src11_valid),               //          .valid
		.in_startofpacket  (cmd_xbar_demux_src11_startofpacket),       //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src11_endofpacket),         //          .endofpacket
		.in_data           (cmd_xbar_demux_src11_data),                //          .data
		.in_channel        (cmd_xbar_demux_src11_channel),             //          .channel
		.out_ready         (agent_pipeline_022_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_022_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_022_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_022_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_022_source0_data),          //          .data
		.out_channel       (agent_pipeline_022_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_023 (
		.clk               (clk_clk),                                                           //       cr0.clk
		.reset             (rst_controller_reset_out_reset),                                    // cr0_reset.reset
		.in_ready          (key_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (key_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (key_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (key_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (key_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_023_source0_ready),                                  //   source0.ready
		.out_valid         (agent_pipeline_023_source0_valid),                                  //          .valid
		.out_startofpacket (agent_pipeline_023_source0_startofpacket),                          //          .startofpacket
		.out_endofpacket   (agent_pipeline_023_source0_endofpacket),                            //          .endofpacket
		.out_data          (agent_pipeline_023_source0_data),                                   //          .data
		.in_empty          (1'b0),                                                              // (terminated)
		.out_empty         (),                                                                  // (terminated)
		.out_error         (),                                                                  // (terminated)
		.in_error          (1'b0),                                                              // (terminated)
		.out_channel       (),                                                                  // (terminated)
		.in_channel        (1'b0)                                                               // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (25),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_024 (
		.clk               (clk_clk),                                  //       cr0.clk
		.reset             (rst_controller_reset_out_reset),           // cr0_reset.reset
		.in_ready          (cmd_xbar_demux_src12_ready),               //     sink0.ready
		.in_valid          (cmd_xbar_demux_src12_valid),               //          .valid
		.in_startofpacket  (cmd_xbar_demux_src12_startofpacket),       //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src12_endofpacket),         //          .endofpacket
		.in_data           (cmd_xbar_demux_src12_data),                //          .data
		.in_channel        (cmd_xbar_demux_src12_channel),             //          .channel
		.out_ready         (agent_pipeline_024_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_024_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_024_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_024_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_024_source0_data),          //          .data
		.out_channel       (agent_pipeline_024_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_025 (
		.clk               (clk_clk),                                                                       //       cr0.clk
		.reset             (rst_controller_reset_out_reset),                                                // cr0_reset.reset
		.in_ready          (signal_selector_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (signal_selector_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (signal_selector_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (signal_selector_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (signal_selector_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_025_source0_ready),                                              //   source0.ready
		.out_valid         (agent_pipeline_025_source0_valid),                                              //          .valid
		.out_startofpacket (agent_pipeline_025_source0_startofpacket),                                      //          .startofpacket
		.out_endofpacket   (agent_pipeline_025_source0_endofpacket),                                        //          .endofpacket
		.out_data          (agent_pipeline_025_source0_data),                                               //          .data
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_channel       (),                                                                              // (terminated)
		.in_channel        (1'b0)                                                                           // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (25),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_026 (
		.clk               (clk_clk),                                  //       cr0.clk
		.reset             (rst_controller_reset_out_reset),           // cr0_reset.reset
		.in_ready          (cmd_xbar_demux_src13_ready),               //     sink0.ready
		.in_valid          (cmd_xbar_demux_src13_valid),               //          .valid
		.in_startofpacket  (cmd_xbar_demux_src13_startofpacket),       //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src13_endofpacket),         //          .endofpacket
		.in_data           (cmd_xbar_demux_src13_data),                //          .data
		.in_channel        (cmd_xbar_demux_src13_channel),             //          .channel
		.out_ready         (agent_pipeline_026_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_026_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_026_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_026_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_026_source0_data),          //          .data
		.out_channel       (agent_pipeline_026_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_027 (
		.clk               (clk_clk),                                                                           //       cr0.clk
		.reset             (rst_controller_reset_out_reset),                                                    // cr0_reset.reset
		.in_ready          (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (modulation_selector_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_027_source0_ready),                                                  //   source0.ready
		.out_valid         (agent_pipeline_027_source0_valid),                                                  //          .valid
		.out_startofpacket (agent_pipeline_027_source0_startofpacket),                                          //          .startofpacket
		.out_endofpacket   (agent_pipeline_027_source0_endofpacket),                                            //          .endofpacket
		.out_data          (agent_pipeline_027_source0_data),                                                   //          .data
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_channel       (),                                                                                  // (terminated)
		.in_channel        (1'b0)                                                                               // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (25),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_028 (
		.clk               (clk_25_in_clk),                            //       cr0.clk
		.reset             (rst_controller_002_reset_out_reset),       // cr0_reset.reset
		.in_ready          (crosser_out_ready),                        //     sink0.ready
		.in_valid          (crosser_out_valid),                        //          .valid
		.in_startofpacket  (crosser_out_startofpacket),                //          .startofpacket
		.in_endofpacket    (crosser_out_endofpacket),                  //          .endofpacket
		.in_data           (crosser_out_data),                         //          .data
		.in_channel        (crosser_out_channel),                      //          .channel
		.out_ready         (agent_pipeline_028_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_028_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_028_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_028_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_028_source0_data),          //          .data
		.out_channel       (agent_pipeline_028_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_029 (
		.clk               (clk_25_in_clk),                                                               //       cr0.clk
		.reset             (rst_controller_002_reset_out_reset),                                          // cr0_reset.reset
		.in_ready          (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (keyboard_keys_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_029_source0_ready),                                            //   source0.ready
		.out_valid         (agent_pipeline_029_source0_valid),                                            //          .valid
		.out_startofpacket (agent_pipeline_029_source0_startofpacket),                                    //          .startofpacket
		.out_endofpacket   (agent_pipeline_029_source0_endofpacket),                                      //          .endofpacket
		.out_data          (agent_pipeline_029_source0_data),                                             //          .data
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_channel       (),                                                                            // (terminated)
		.in_channel        (1'b0)                                                                         // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (25),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_030 (
		.clk               (clk_40_in_clk),                            //       cr0.clk
		.reset             (rst_controller_003_reset_out_reset),       // cr0_reset.reset
		.in_ready          (crosser_001_out_ready),                    //     sink0.ready
		.in_valid          (crosser_001_out_valid),                    //          .valid
		.in_startofpacket  (crosser_001_out_startofpacket),            //          .startofpacket
		.in_endofpacket    (crosser_001_out_endofpacket),              //          .endofpacket
		.in_data           (crosser_001_out_data),                     //          .data
		.in_channel        (crosser_001_out_channel),                  //          .channel
		.out_ready         (agent_pipeline_030_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_030_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_030_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_030_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_030_source0_data),          //          .data
		.out_channel       (agent_pipeline_030_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_031 (
		.clk               (clk_40_in_clk),                                                           //       cr0.clk
		.reset             (rst_controller_003_reset_out_reset),                                      // cr0_reset.reset
		.in_ready          (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (mouse_pos_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_031_source0_ready),                                        //   source0.ready
		.out_valid         (agent_pipeline_031_source0_valid),                                        //          .valid
		.out_startofpacket (agent_pipeline_031_source0_startofpacket),                                //          .startofpacket
		.out_endofpacket   (agent_pipeline_031_source0_endofpacket),                                  //          .endofpacket
		.out_data          (agent_pipeline_031_source0_data),                                         //          .data
		.in_empty          (1'b0),                                                                    // (terminated)
		.out_empty         (),                                                                        // (terminated)
		.out_error         (),                                                                        // (terminated)
		.in_error          (1'b0),                                                                    // (terminated)
		.out_channel       (),                                                                        // (terminated)
		.in_channel        (1'b0)                                                                     // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (25),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_032 (
		.clk               (clk_clk),                                  //       cr0.clk
		.reset             (rst_controller_reset_out_reset),           // cr0_reset.reset
		.in_ready          (cmd_xbar_demux_src16_ready),               //     sink0.ready
		.in_valid          (cmd_xbar_demux_src16_valid),               //          .valid
		.in_startofpacket  (cmd_xbar_demux_src16_startofpacket),       //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src16_endofpacket),         //          .endofpacket
		.in_data           (cmd_xbar_demux_src16_data),                //          .data
		.in_channel        (cmd_xbar_demux_src16_channel),             //          .channel
		.out_ready         (agent_pipeline_032_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_032_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_032_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_032_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_032_source0_data),          //          .data
		.out_channel       (agent_pipeline_032_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_033 (
		.clk               (clk_clk),                                                                //       cr0.clk
		.reset             (rst_controller_reset_out_reset),                                         // cr0_reset.reset
		.in_ready          (div_freq_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (div_freq_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (div_freq_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (div_freq_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (div_freq_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_033_source0_ready),                                       //   source0.ready
		.out_valid         (agent_pipeline_033_source0_valid),                                       //          .valid
		.out_startofpacket (agent_pipeline_033_source0_startofpacket),                               //          .startofpacket
		.out_endofpacket   (agent_pipeline_033_source0_endofpacket),                                 //          .endofpacket
		.out_data          (agent_pipeline_033_source0_data),                                        //          .data
		.in_empty          (1'b0),                                                                   // (terminated)
		.out_empty         (),                                                                       // (terminated)
		.out_error         (),                                                                       // (terminated)
		.in_error          (1'b0),                                                                   // (terminated)
		.out_channel       (),                                                                       // (terminated)
		.in_channel        (1'b0)                                                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (25),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_034 (
		.clk               (clk_clk),                                  //       cr0.clk
		.reset             (rst_controller_reset_out_reset),           // cr0_reset.reset
		.in_ready          (cmd_xbar_demux_src17_ready),               //     sink0.ready
		.in_valid          (cmd_xbar_demux_src17_valid),               //          .valid
		.in_startofpacket  (cmd_xbar_demux_src17_startofpacket),       //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src17_endofpacket),         //          .endofpacket
		.in_data           (cmd_xbar_demux_src17_data),                //          .data
		.in_channel        (cmd_xbar_demux_src17_channel),             //          .channel
		.out_ready         (agent_pipeline_034_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_034_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_034_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_034_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_034_source0_data),          //          .data
		.out_channel       (agent_pipeline_034_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_035 (
		.clk               (clk_clk),                                                                 //       cr0.clk
		.reset             (rst_controller_reset_out_reset),                                          // cr0_reset.reset
		.in_ready          (audio_sel_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (audio_sel_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (audio_sel_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (audio_sel_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (audio_sel_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_035_source0_ready),                                        //   source0.ready
		.out_valid         (agent_pipeline_035_source0_valid),                                        //          .valid
		.out_startofpacket (agent_pipeline_035_source0_startofpacket),                                //          .startofpacket
		.out_endofpacket   (agent_pipeline_035_source0_endofpacket),                                  //          .endofpacket
		.out_data          (agent_pipeline_035_source0_data),                                         //          .data
		.in_empty          (1'b0),                                                                    // (terminated)
		.out_empty         (),                                                                        // (terminated)
		.out_error         (),                                                                        // (terminated)
		.in_error          (1'b0),                                                                    // (terminated)
		.out_channel       (),                                                                        // (terminated)
		.in_channel        (1'b0)                                                                     // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (25),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_036 (
		.clk               (cpu_clk_for_sdram_clk),                    //       cr0.clk
		.reset             (rst_controller_004_reset_out_reset),       // cr0_reset.reset
		.in_ready          (crosser_002_out_ready),                    //     sink0.ready
		.in_valid          (crosser_002_out_valid),                    //          .valid
		.in_startofpacket  (crosser_002_out_startofpacket),            //          .startofpacket
		.in_endofpacket    (crosser_002_out_endofpacket),              //          .endofpacket
		.in_data           (crosser_002_out_data),                     //          .data
		.in_channel        (crosser_002_out_channel),                  //          .channel
		.out_ready         (agent_pipeline_036_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_036_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_036_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_036_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_036_source0_data),          //          .data
		.out_channel       (agent_pipeline_036_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_037 (
		.clk               (cpu_clk_for_sdram_clk),                                                               //       cr0.clk
		.reset             (rst_controller_004_reset_out_reset),                                                  // cr0_reset.reset
		.in_ready          (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (vga_to_nios_2_datamaster_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_037_source0_ready),                                                    //   source0.ready
		.out_valid         (agent_pipeline_037_source0_valid),                                                    //          .valid
		.out_startofpacket (agent_pipeline_037_source0_startofpacket),                                            //          .startofpacket
		.out_endofpacket   (agent_pipeline_037_source0_endofpacket),                                              //          .endofpacket
		.out_data          (agent_pipeline_037_source0_data),                                                     //          .data
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_channel       (),                                                                                    // (terminated)
		.in_channel        (1'b0)                                                                                 // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (25),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_038 (
		.clk               (clk_clk),                                  //       cr0.clk
		.reset             (rst_controller_reset_out_reset),           // cr0_reset.reset
		.in_ready          (cmd_xbar_demux_src19_ready),               //     sink0.ready
		.in_valid          (cmd_xbar_demux_src19_valid),               //          .valid
		.in_startofpacket  (cmd_xbar_demux_src19_startofpacket),       //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src19_endofpacket),         //          .endofpacket
		.in_data           (cmd_xbar_demux_src19_data),                //          .data
		.in_channel        (cmd_xbar_demux_src19_channel),             //          .channel
		.out_ready         (agent_pipeline_038_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_038_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_038_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_038_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_038_source0_data),          //          .data
		.out_channel       (agent_pipeline_038_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_039 (
		.clk               (clk_clk),                                                                   //       cr0.clk
		.reset             (rst_controller_reset_out_reset),                                            // cr0_reset.reset
		.in_ready          (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (audio_wrclk_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_039_source0_ready),                                          //   source0.ready
		.out_valid         (agent_pipeline_039_source0_valid),                                          //          .valid
		.out_startofpacket (agent_pipeline_039_source0_startofpacket),                                  //          .startofpacket
		.out_endofpacket   (agent_pipeline_039_source0_endofpacket),                                    //          .endofpacket
		.out_data          (agent_pipeline_039_source0_data),                                           //          .data
		.in_empty          (1'b0),                                                                      // (terminated)
		.out_empty         (),                                                                          // (terminated)
		.out_error         (),                                                                          // (terminated)
		.in_error          (1'b0),                                                                      // (terminated)
		.out_channel       (),                                                                          // (terminated)
		.in_channel        (1'b0)                                                                       // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (25),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_040 (
		.clk               (clk_clk),                                  //       cr0.clk
		.reset             (rst_controller_reset_out_reset),           // cr0_reset.reset
		.in_ready          (cmd_xbar_demux_src20_ready),               //     sink0.ready
		.in_valid          (cmd_xbar_demux_src20_valid),               //          .valid
		.in_startofpacket  (cmd_xbar_demux_src20_startofpacket),       //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src20_endofpacket),         //          .endofpacket
		.in_data           (cmd_xbar_demux_src20_data),                //          .data
		.in_channel        (cmd_xbar_demux_src20_channel),             //          .channel
		.out_ready         (agent_pipeline_040_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_040_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_040_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_040_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_040_source0_data),          //          .data
		.out_channel       (agent_pipeline_040_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_041 (
		.clk               (clk_clk),                                                                   //       cr0.clk
		.reset             (rst_controller_reset_out_reset),                                            // cr0_reset.reset
		.in_ready          (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (audio_wrreq_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_041_source0_ready),                                          //   source0.ready
		.out_valid         (agent_pipeline_041_source0_valid),                                          //          .valid
		.out_startofpacket (agent_pipeline_041_source0_startofpacket),                                  //          .startofpacket
		.out_endofpacket   (agent_pipeline_041_source0_endofpacket),                                    //          .endofpacket
		.out_data          (agent_pipeline_041_source0_data),                                           //          .data
		.in_empty          (1'b0),                                                                      // (terminated)
		.out_empty         (),                                                                          // (terminated)
		.out_error         (),                                                                          // (terminated)
		.in_error          (1'b0),                                                                      // (terminated)
		.out_channel       (),                                                                          // (terminated)
		.in_channel        (1'b0)                                                                       // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (96),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (25),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_042 (
		.clk               (cpu_clk_for_sdram_clk),                    //       cr0.clk
		.reset             (rst_controller_004_reset_out_reset),       // cr0_reset.reset
		.in_ready          (burst_adapter_source0_ready),              //     sink0.ready
		.in_valid          (burst_adapter_source0_valid),              //          .valid
		.in_startofpacket  (burst_adapter_source0_startofpacket),      //          .startofpacket
		.in_endofpacket    (burst_adapter_source0_endofpacket),        //          .endofpacket
		.in_data           (burst_adapter_source0_data),               //          .data
		.in_channel        (burst_adapter_source0_channel),            //          .channel
		.out_ready         (agent_pipeline_042_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_042_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_042_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_042_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_042_source0_data),          //          .data
		.out_channel       (agent_pipeline_042_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (96),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_043 (
		.clk               (cpu_clk_for_sdram_clk),                                               //       cr0.clk
		.reset             (rst_controller_004_reset_out_reset),                                  // cr0_reset.reset
		.in_ready          (sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_043_source0_ready),                                    //   source0.ready
		.out_valid         (agent_pipeline_043_source0_valid),                                    //          .valid
		.out_startofpacket (agent_pipeline_043_source0_startofpacket),                            //          .startofpacket
		.out_endofpacket   (agent_pipeline_043_source0_endofpacket),                              //          .endofpacket
		.out_data          (agent_pipeline_043_source0_data),                                     //          .data
		.in_empty          (1'b0),                                                                // (terminated)
		.out_empty         (),                                                                    // (terminated)
		.out_error         (),                                                                    // (terminated)
		.in_error          (1'b0),                                                                // (terminated)
		.out_channel       (),                                                                    // (terminated)
		.in_channel        (1'b0)                                                                 // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (25),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_044 (
		.clk               (clk_clk),                                  //       cr0.clk
		.reset             (rst_controller_reset_out_reset),           // cr0_reset.reset
		.in_ready          (cmd_xbar_demux_src22_ready),               //     sink0.ready
		.in_valid          (cmd_xbar_demux_src22_valid),               //          .valid
		.in_startofpacket  (cmd_xbar_demux_src22_startofpacket),       //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src22_endofpacket),         //          .endofpacket
		.in_data           (cmd_xbar_demux_src22_data),                //          .data
		.in_channel        (cmd_xbar_demux_src22_channel),             //          .channel
		.out_ready         (agent_pipeline_044_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_044_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_044_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_044_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_044_source0_data),          //          .data
		.out_channel       (agent_pipeline_044_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_045 (
		.clk               (clk_clk),                                                                              //       cr0.clk
		.reset             (rst_controller_reset_out_reset),                                                       // cr0_reset.reset
		.in_ready          (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (lfsr_clk_interrupt_gen_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_045_source0_ready),                                                     //   source0.ready
		.out_valid         (agent_pipeline_045_source0_valid),                                                     //          .valid
		.out_startofpacket (agent_pipeline_045_source0_startofpacket),                                             //          .startofpacket
		.out_endofpacket   (agent_pipeline_045_source0_endofpacket),                                               //          .endofpacket
		.out_data          (agent_pipeline_045_source0_data),                                                      //          .data
		.in_empty          (1'b0),                                                                                 // (terminated)
		.out_empty         (),                                                                                     // (terminated)
		.out_error         (),                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                 // (terminated)
		.out_channel       (),                                                                                     // (terminated)
		.in_channel        (1'b0)                                                                                  // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (25),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_046 (
		.clk               (clk_clk),                                  //       cr0.clk
		.reset             (rst_controller_reset_out_reset),           // cr0_reset.reset
		.in_ready          (cmd_xbar_demux_src23_ready),               //     sink0.ready
		.in_valid          (cmd_xbar_demux_src23_valid),               //          .valid
		.in_startofpacket  (cmd_xbar_demux_src23_startofpacket),       //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src23_endofpacket),         //          .endofpacket
		.in_data           (cmd_xbar_demux_src23_data),                //          .data
		.in_channel        (cmd_xbar_demux_src23_channel),             //          .channel
		.out_ready         (agent_pipeline_046_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_046_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_046_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_046_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_046_source0_data),          //          .data
		.out_channel       (agent_pipeline_046_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_047 (
		.clk               (clk_clk),                                                                //       cr0.clk
		.reset             (rst_controller_reset_out_reset),                                         // cr0_reset.reset
		.in_ready          (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (lfsr_val_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_047_source0_ready),                                       //   source0.ready
		.out_valid         (agent_pipeline_047_source0_valid),                                       //          .valid
		.out_startofpacket (agent_pipeline_047_source0_startofpacket),                               //          .startofpacket
		.out_endofpacket   (agent_pipeline_047_source0_endofpacket),                                 //          .endofpacket
		.out_data          (agent_pipeline_047_source0_data),                                        //          .data
		.in_empty          (1'b0),                                                                   // (terminated)
		.out_empty         (),                                                                       // (terminated)
		.out_error         (),                                                                       // (terminated)
		.in_error          (1'b0),                                                                   // (terminated)
		.out_channel       (),                                                                       // (terminated)
		.in_channel        (1'b0)                                                                    // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (25),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_048 (
		.clk               (clk_clk),                                  //       cr0.clk
		.reset             (rst_controller_reset_out_reset),           // cr0_reset.reset
		.in_ready          (cmd_xbar_demux_src24_ready),               //     sink0.ready
		.in_valid          (cmd_xbar_demux_src24_valid),               //          .valid
		.in_startofpacket  (cmd_xbar_demux_src24_startofpacket),       //          .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src24_endofpacket),         //          .endofpacket
		.in_data           (cmd_xbar_demux_src24_data),                //          .data
		.in_channel        (cmd_xbar_demux_src24_channel),             //          .channel
		.out_ready         (agent_pipeline_048_source0_ready),         //   source0.ready
		.out_valid         (agent_pipeline_048_source0_valid),         //          .valid
		.out_startofpacket (agent_pipeline_048_source0_startofpacket), //          .startofpacket
		.out_endofpacket   (agent_pipeline_048_source0_endofpacket),   //          .endofpacket
		.out_data          (agent_pipeline_048_source0_data),          //          .data
		.out_channel       (agent_pipeline_048_source0_channel),       //          .channel
		.in_empty          (1'b0),                                     // (terminated)
		.out_empty         (),                                         // (terminated)
		.out_error         (),                                         // (terminated)
		.in_error          (1'b0)                                      // (terminated)
	);

	altera_avalon_st_pipeline_stage #(
		.SYMBOLS_PER_BEAT (1),
		.BITS_PER_SYMBOL  (114),
		.USE_PACKETS      (1),
		.USE_EMPTY        (0),
		.EMPTY_WIDTH      (0),
		.CHANNEL_WIDTH    (0),
		.PACKET_WIDTH     (2),
		.ERROR_WIDTH      (0),
		.PIPELINE_READY   (1)
	) agent_pipeline_049 (
		.clk               (clk_clk),                                                                     //       cr0.clk
		.reset             (rst_controller_reset_out_reset),                                              // cr0_reset.reset
		.in_ready          (dds_increment_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //     sink0.ready
		.in_valid          (dds_increment_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.in_startofpacket  (dds_increment_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.in_endofpacket    (dds_increment_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.in_data           (dds_increment_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.out_ready         (agent_pipeline_049_source0_ready),                                            //   source0.ready
		.out_valid         (agent_pipeline_049_source0_valid),                                            //          .valid
		.out_startofpacket (agent_pipeline_049_source0_startofpacket),                                    //          .startofpacket
		.out_endofpacket   (agent_pipeline_049_source0_endofpacket),                                      //          .endofpacket
		.out_data          (agent_pipeline_049_source0_data),                                             //          .data
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_channel       (),                                                                            // (terminated)
		.in_channel        (1'b0)                                                                         // (terminated)
	);

	DE2_QSYS_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.sender_irq    (cpu_d_irq_irq)                       //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (cpu_clk_for_sdram_clk),              //       receiver_clk.clk
		.sender_clk     (clk_clk),                            //         sender_clk.clk
		.receiver_reset (~reset_reset_n),                     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	assign vga_vga_clk_clk = clk_40_in_clk;

endmodule
